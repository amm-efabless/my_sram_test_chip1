// This is the unpowered netlist.
module wishbone_sram (sram_selected,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 output sram_selected;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \ram_controller.DO[0] ;
 wire \ram_controller.DO[10] ;
 wire \ram_controller.DO[11] ;
 wire \ram_controller.DO[12] ;
 wire \ram_controller.DO[13] ;
 wire \ram_controller.DO[14] ;
 wire \ram_controller.DO[15] ;
 wire \ram_controller.DO[16] ;
 wire \ram_controller.DO[17] ;
 wire \ram_controller.DO[18] ;
 wire \ram_controller.DO[19] ;
 wire \ram_controller.DO[1] ;
 wire \ram_controller.DO[20] ;
 wire \ram_controller.DO[21] ;
 wire \ram_controller.DO[22] ;
 wire \ram_controller.DO[23] ;
 wire \ram_controller.DO[24] ;
 wire \ram_controller.DO[25] ;
 wire \ram_controller.DO[26] ;
 wire \ram_controller.DO[27] ;
 wire \ram_controller.DO[28] ;
 wire \ram_controller.DO[29] ;
 wire \ram_controller.DO[2] ;
 wire \ram_controller.DO[30] ;
 wire \ram_controller.DO[31] ;
 wire \ram_controller.DO[3] ;
 wire \ram_controller.DO[4] ;
 wire \ram_controller.DO[5] ;
 wire \ram_controller.DO[6] ;
 wire \ram_controller.DO[7] ;
 wire \ram_controller.DO[8] ;
 wire \ram_controller.DO[9] ;
 wire \ram_controller.EN ;
 wire \ram_controller.R_WB ;
 wire \ram_controller.wbs_ack_o ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_800 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_2_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_2_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_2_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_2_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Right_164 ();
 EFSRAM_1024x32_wrapper SRAM_0 (.WLBI(net92),
    .WLOFF(net93),
    .CLKin(clknet_1_1__leaf_wb_clk_i),
    .EN(\ram_controller.EN ),
    .R_WB(\ram_controller.R_WB ),
    .SM(net87),
    .TM(net91),
    .ScanInDR(net90),
    .ScanInDL(net89),
    .ScanInCC(net88),
    .vpwrpc(net95),
    .vpwrac(net94),
    .AD({net155,
    net163,
    net165,
    net167,
    net169,
    net171,
    net173,
    net175,
    net177,
    net179}),
    .BEN({net190,
    net190,
    net190,
    net190,
    net190,
    net190,
    net190,
    net190,
    net187,
    net187,
    net187,
    net187,
    net187,
    net187,
    net187,
    net187,
    net181,
    net181,
    net181,
    net181,
    net181,
    net181,
    net181,
    net181,
    net184,
    net184,
    net184,
    net184,
    net184,
    net184,
    net184,
    net184}),
    .DI({net129,
    net125,
    net119,
    net111,
    net107,
    net101,
    net161,
    net157,
    net151,
    net153,
    net149,
    net147,
    net139,
    net141,
    net143,
    net145,
    net99,
    net113,
    net123,
    net131,
    net97,
    net109,
    net121,
    net127,
    net133,
    net135,
    net137,
    net159,
    net103,
    net105,
    net115,
    net117}),
    .DO({\ram_controller.DO[31] ,
    \ram_controller.DO[30] ,
    \ram_controller.DO[29] ,
    \ram_controller.DO[28] ,
    \ram_controller.DO[27] ,
    \ram_controller.DO[26] ,
    \ram_controller.DO[25] ,
    \ram_controller.DO[24] ,
    \ram_controller.DO[23] ,
    \ram_controller.DO[22] ,
    \ram_controller.DO[21] ,
    \ram_controller.DO[20] ,
    \ram_controller.DO[19] ,
    \ram_controller.DO[18] ,
    \ram_controller.DO[17] ,
    \ram_controller.DO[16] ,
    \ram_controller.DO[15] ,
    \ram_controller.DO[14] ,
    \ram_controller.DO[13] ,
    \ram_controller.DO[12] ,
    \ram_controller.DO[11] ,
    \ram_controller.DO[10] ,
    \ram_controller.DO[9] ,
    \ram_controller.DO[8] ,
    \ram_controller.DO[7] ,
    \ram_controller.DO[6] ,
    \ram_controller.DO[5] ,
    \ram_controller.DO[4] ,
    \ram_controller.DO[3] ,
    \ram_controller.DO[2] ,
    \ram_controller.DO[1] ,
    \ram_controller.DO[0] }));
 sky130_fd_sc_hd__conb_1 SRAM_0_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 SRAM_0_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 SRAM_0_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 SRAM_0_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 SRAM_0_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 SRAM_0_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 SRAM_0_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 SRAM_0_94 (.HI(net94));
 sky130_fd_sc_hd__conb_1 SRAM_0_95 (.HI(net95));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_2_687 ();
 sky130_fd_sc_hd__nor2b_4 _049_ (.A(net193),
    .B_N(net4),
    .Y(_028_));
 sky130_fd_sc_hd__clkbuf_4 _050_ (.A(_028_),
    .X(net53));
 sky130_fd_sc_hd__and2_1 _051_ (.A(\ram_controller.DO[0] ),
    .B(net53),
    .X(_029_));
 sky130_fd_sc_hd__buf_1 _052_ (.A(_029_),
    .X(net55));
 sky130_fd_sc_hd__and2_1 _053_ (.A(\ram_controller.DO[1] ),
    .B(net53),
    .X(_030_));
 sky130_fd_sc_hd__buf_1 _054_ (.A(_030_),
    .X(net66));
 sky130_fd_sc_hd__and2_1 _055_ (.A(\ram_controller.DO[2] ),
    .B(net53),
    .X(_031_));
 sky130_fd_sc_hd__buf_1 _056_ (.A(_031_),
    .X(net77));
 sky130_fd_sc_hd__and2_1 _057_ (.A(\ram_controller.DO[3] ),
    .B(net53),
    .X(_032_));
 sky130_fd_sc_hd__buf_1 _058_ (.A(_032_),
    .X(net80));
 sky130_fd_sc_hd__and2_1 _059_ (.A(\ram_controller.DO[4] ),
    .B(net53),
    .X(_033_));
 sky130_fd_sc_hd__buf_1 _060_ (.A(_033_),
    .X(net81));
 sky130_fd_sc_hd__and2_1 _061_ (.A(\ram_controller.DO[5] ),
    .B(net53),
    .X(_034_));
 sky130_fd_sc_hd__buf_1 _062_ (.A(_034_),
    .X(net82));
 sky130_fd_sc_hd__and2_1 _063_ (.A(\ram_controller.DO[6] ),
    .B(net53),
    .X(_035_));
 sky130_fd_sc_hd__buf_1 _064_ (.A(_035_),
    .X(net83));
 sky130_fd_sc_hd__and2_1 _065_ (.A(\ram_controller.DO[7] ),
    .B(net53),
    .X(_036_));
 sky130_fd_sc_hd__buf_1 _066_ (.A(_036_),
    .X(net84));
 sky130_fd_sc_hd__and2_1 _067_ (.A(\ram_controller.DO[8] ),
    .B(net53),
    .X(_037_));
 sky130_fd_sc_hd__buf_1 _068_ (.A(_037_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 _069_ (.A(_028_),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _070_ (.A(\ram_controller.DO[9] ),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__buf_1 _071_ (.A(_039_),
    .X(net86));
 sky130_fd_sc_hd__and2_1 _072_ (.A(\ram_controller.DO[10] ),
    .B(_038_),
    .X(_002_));
 sky130_fd_sc_hd__buf_1 _073_ (.A(_002_),
    .X(net56));
 sky130_fd_sc_hd__and2_1 _074_ (.A(\ram_controller.DO[11] ),
    .B(_038_),
    .X(_003_));
 sky130_fd_sc_hd__buf_1 _075_ (.A(_003_),
    .X(net57));
 sky130_fd_sc_hd__and2_1 _076_ (.A(\ram_controller.DO[12] ),
    .B(_038_),
    .X(_004_));
 sky130_fd_sc_hd__buf_1 _077_ (.A(_004_),
    .X(net58));
 sky130_fd_sc_hd__and2_1 _078_ (.A(\ram_controller.DO[13] ),
    .B(_038_),
    .X(_005_));
 sky130_fd_sc_hd__buf_1 _079_ (.A(_005_),
    .X(net59));
 sky130_fd_sc_hd__and2_1 _080_ (.A(\ram_controller.DO[14] ),
    .B(_038_),
    .X(_006_));
 sky130_fd_sc_hd__buf_1 _081_ (.A(_006_),
    .X(net60));
 sky130_fd_sc_hd__and2_1 _082_ (.A(\ram_controller.DO[15] ),
    .B(_038_),
    .X(_007_));
 sky130_fd_sc_hd__buf_1 _083_ (.A(_007_),
    .X(net61));
 sky130_fd_sc_hd__and2_1 _084_ (.A(\ram_controller.DO[16] ),
    .B(_038_),
    .X(_008_));
 sky130_fd_sc_hd__buf_1 _085_ (.A(_008_),
    .X(net62));
 sky130_fd_sc_hd__and2_1 _086_ (.A(\ram_controller.DO[17] ),
    .B(_038_),
    .X(_009_));
 sky130_fd_sc_hd__buf_1 _087_ (.A(_009_),
    .X(net63));
 sky130_fd_sc_hd__and2_1 _088_ (.A(\ram_controller.DO[18] ),
    .B(_038_),
    .X(_010_));
 sky130_fd_sc_hd__buf_1 _089_ (.A(_010_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 _090_ (.A(_028_),
    .X(_011_));
 sky130_fd_sc_hd__and2_1 _091_ (.A(\ram_controller.DO[19] ),
    .B(_011_),
    .X(_012_));
 sky130_fd_sc_hd__buf_1 _092_ (.A(_012_),
    .X(net65));
 sky130_fd_sc_hd__and2_1 _093_ (.A(\ram_controller.DO[20] ),
    .B(_011_),
    .X(_013_));
 sky130_fd_sc_hd__buf_1 _094_ (.A(_013_),
    .X(net67));
 sky130_fd_sc_hd__and2_1 _095_ (.A(\ram_controller.DO[21] ),
    .B(_011_),
    .X(_014_));
 sky130_fd_sc_hd__buf_1 _096_ (.A(_014_),
    .X(net68));
 sky130_fd_sc_hd__and2_1 _097_ (.A(\ram_controller.DO[22] ),
    .B(_011_),
    .X(_015_));
 sky130_fd_sc_hd__buf_1 _098_ (.A(_015_),
    .X(net69));
 sky130_fd_sc_hd__and2_1 _099_ (.A(\ram_controller.DO[23] ),
    .B(_011_),
    .X(_016_));
 sky130_fd_sc_hd__buf_1 _100_ (.A(_016_),
    .X(net70));
 sky130_fd_sc_hd__and2_1 _101_ (.A(\ram_controller.DO[24] ),
    .B(_011_),
    .X(_017_));
 sky130_fd_sc_hd__buf_1 _102_ (.A(_017_),
    .X(net71));
 sky130_fd_sc_hd__and2_1 _103_ (.A(\ram_controller.DO[25] ),
    .B(_011_),
    .X(_018_));
 sky130_fd_sc_hd__buf_1 _104_ (.A(_018_),
    .X(net72));
 sky130_fd_sc_hd__and2_1 _105_ (.A(\ram_controller.DO[26] ),
    .B(_011_),
    .X(_019_));
 sky130_fd_sc_hd__buf_1 _106_ (.A(_019_),
    .X(net73));
 sky130_fd_sc_hd__and2_1 _107_ (.A(\ram_controller.DO[27] ),
    .B(_011_),
    .X(_020_));
 sky130_fd_sc_hd__buf_1 _108_ (.A(_020_),
    .X(net74));
 sky130_fd_sc_hd__and2_1 _109_ (.A(\ram_controller.DO[28] ),
    .B(_011_),
    .X(_021_));
 sky130_fd_sc_hd__buf_1 _110_ (.A(_021_),
    .X(net75));
 sky130_fd_sc_hd__and2_1 _111_ (.A(\ram_controller.DO[29] ),
    .B(_028_),
    .X(_022_));
 sky130_fd_sc_hd__buf_1 _112_ (.A(_022_),
    .X(net76));
 sky130_fd_sc_hd__and2_1 _113_ (.A(\ram_controller.DO[30] ),
    .B(_028_),
    .X(_023_));
 sky130_fd_sc_hd__buf_1 _114_ (.A(_023_),
    .X(net78));
 sky130_fd_sc_hd__and2_1 _115_ (.A(\ram_controller.DO[31] ),
    .B(_028_),
    .X(_024_));
 sky130_fd_sc_hd__buf_1 _116_ (.A(_024_),
    .X(net79));
 sky130_fd_sc_hd__clkinv_4 _117_ (.A(net52),
    .Y(\ram_controller.R_WB ));
 sky130_fd_sc_hd__and2_1 _118_ (.A(\ram_controller.wbs_ack_o ),
    .B(_028_),
    .X(_025_));
 sky130_fd_sc_hd__buf_1 _119_ (.A(_025_),
    .X(net54));
 sky130_fd_sc_hd__and3_1 _120_ (.A(net14),
    .B(net51),
    .C(net194),
    .X(_026_));
 sky130_fd_sc_hd__buf_4 _121_ (.A(net195),
    .X(\ram_controller.EN ));
 sky130_fd_sc_hd__and4b_1 _122_ (.A_N(\ram_controller.wbs_ack_o ),
    .B(net14),
    .C(net51),
    .D(net194),
    .X(_027_));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(_027_),
    .X(_000_));
 sky130_fd_sc_hd__inv_2 _124_ (.A(net1),
    .Y(_001_));
 sky130_fd_sc_hd__dfrtp_1 _125_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_000_),
    .RESET_B(_001_),
    .Q(\ram_controller.wbs_ack_o ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net201),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net37),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_026_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(wbs_we_i),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(wbs_dat_i[15]),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(wbs_dat_i[14]),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(wbs_dat_i[13]),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(wbs_dat_i[12]),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(wbs_dat_i[11]),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(wbs_dat_i[10]),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(wbs_dat_i[9]),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(wbs_dat_i[8]),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net222),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(wbs_dat_i[7]),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(wbs_dat_i[6]),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(wbs_dat_i[19]),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(wbs_dat_i[18]),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(wbs_dat_i[5]),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(wbs_dat_i[17]),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(wbs_dat_i[16]),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(wbs_dat_i[20]),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(wbs_dat_i[3]),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(wbs_dat_i[23]),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net34),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(wbs_dat_i[21]),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(wbs_dat_i[26]),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(wbs_dat_i[22]),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(wbs_dat_i[4]),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(wbs_dat_i[24]),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(wbs_dat_i[2]),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(wbs_dat_i[25]),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(wbs_dat_i[27]),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(wbs_dat_i[28]),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(wbs_dat_i[1]),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net202),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(wbs_dat_i[0]),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(wbs_dat_i[29]),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(wbs_dat_i[30]),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(wbs_dat_i[31]),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(wbs_adr_i[9]),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(wbs_adr_i[8]),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(wbs_adr_i[7]),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(wbs_adr_i[6]),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(wbs_adr_i[5]),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(wbs_adr_i[4]),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net16),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(wbs_adr_i[3]),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(wbs_adr_i[2]),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(wbs_adr_i[1]),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(wbs_adr_i[0]),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net223),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net35),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net198),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net20),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net224),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net17),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net26),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net225),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net15),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net226),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net36),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net203),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net46),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net199),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net19),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net227),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net197),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net38),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net204),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net45),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net228),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net39),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net200),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net18),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net205),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net44),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net206),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net21),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net43),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net209),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net42),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net207),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net25),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net208),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net24),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net210),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net23),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net211),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net216),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net22),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net212),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net27),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net215),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net28),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net214),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net30),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net217),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net29),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net229),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net33),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net13),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net219),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net31),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net218),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net41),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net221),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net32),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net230),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net12),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net231),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net213),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net11),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net232),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net10),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net233),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net9),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net234),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net8),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net235),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net7),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net236),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net40),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net6),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net237),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net5),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net238),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net2),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_12 hold86 (.A(net48),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(wbs_sel_i[1]),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__buf_12 hold89 (.A(net47),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net220),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(wbs_sel_i[0]),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__buf_12 hold92 (.A(net49),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(wbs_sel_i[2]),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__buf_12 hold95 (.A(net50),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(wbs_sel_i[3]),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(wbs_adr_i[14]),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net3),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_028_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(net166),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(net164),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(net162),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(net154),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(wbs_cyc_i),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(net116),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(net108),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(net96),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(net130),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(net122),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(net178),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(net112),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(net98),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(net144),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(net142),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(net140),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(net138),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(net114),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(net146),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(net148),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(net152),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(net192),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(net150),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(net156),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(net160),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(net100),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(net106),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(net110),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(net118),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(net104),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(net124),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(net128),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(wbs_adr_i[15]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input40 (.A(net102),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(net158),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(net136),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(net134),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(net132),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(net126),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(net120),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(net183),
    .X(net47));
 sky130_fd_sc_hd__buf_12 input48 (.A(net180),
    .X(net48));
 sky130_fd_sc_hd__buf_12 input49 (.A(net186),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(net176),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input50 (.A(net189),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(wbs_stb_i),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(net196),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input6 (.A(net174),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(net172),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(net170),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(net168),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(sram_selected));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(wbs_dat_o[9]));
endmodule

