magic
tech sky130A
magscale 1 2
timestamp 1715241548
<< viali >>
rect 65625 52445 65659 52479
rect 65901 52445 65935 52479
rect 65625 50269 65659 50303
rect 65625 49589 65659 49623
rect 65625 49181 65659 49215
rect 65625 47005 65659 47039
rect 65901 46937 65935 46971
rect 65625 43741 65659 43775
rect 68017 42721 68051 42755
rect 65625 42653 65659 42687
rect 68661 42653 68695 42687
rect 67097 41769 67131 41803
rect 67741 41565 67775 41599
rect 66453 40681 66487 40715
rect 67097 40477 67131 40511
rect 65625 39593 65659 39627
rect 66269 39389 66303 39423
rect 65625 38505 65659 38539
rect 66269 38301 66303 38335
rect 66269 37213 66303 37247
rect 65625 37145 65659 37179
rect 65625 36329 65659 36363
rect 66269 36125 66303 36159
rect 66545 35717 66579 35751
rect 65809 35649 65843 35683
rect 65625 35241 65659 35275
rect 66269 35037 66303 35071
rect 66913 34153 66947 34187
rect 65625 33881 65659 33915
rect 65625 33609 65659 33643
rect 66269 33405 66303 33439
rect 65625 33065 65659 33099
rect 66269 32861 66303 32895
rect 65625 31977 65659 32011
rect 66269 31773 66303 31807
rect 65625 30889 65659 30923
rect 66269 30685 66303 30719
rect 65625 29801 65659 29835
rect 66269 29597 66303 29631
rect 65625 28713 65659 28747
rect 66269 28509 66303 28543
rect 65625 27557 65659 27591
rect 66269 27421 66303 27455
rect 66637 27013 66671 27047
rect 65809 26945 65843 26979
rect 65625 26537 65659 26571
rect 66269 26333 66303 26367
rect 65625 24361 65659 24395
rect 66269 24157 66303 24191
rect 65625 23817 65659 23851
rect 66269 23613 66303 23647
rect 65625 23273 65659 23307
rect 66269 23069 66303 23103
rect 23673 5865 23707 5899
rect 26157 5865 26191 5899
rect 48145 5865 48179 5899
rect 48881 5865 48915 5899
rect 51089 5865 51123 5899
rect 54033 5865 54067 5899
rect 23305 5729 23339 5763
rect 23765 5729 23799 5763
rect 24317 5729 24351 5763
rect 24777 5729 24811 5763
rect 44925 5729 44959 5763
rect 48973 5729 49007 5763
rect 55229 5729 55263 5763
rect 56517 5729 56551 5763
rect 57805 5729 57839 5763
rect 58173 5729 58207 5763
rect 59369 5729 59403 5763
rect 61669 5729 61703 5763
rect 65073 5729 65107 5763
rect 66177 5729 66211 5763
rect 68477 5729 68511 5763
rect 23489 5661 23523 5695
rect 23949 5661 23983 5695
rect 24501 5661 24535 5695
rect 24961 5661 24995 5695
rect 25881 5661 25915 5695
rect 25973 5661 26007 5695
rect 40417 5661 40451 5695
rect 42349 5661 42383 5695
rect 43545 5661 43579 5695
rect 43821 5661 43855 5695
rect 44465 5661 44499 5695
rect 45569 5661 45603 5695
rect 45661 5661 45695 5695
rect 46397 5661 46431 5695
rect 47041 5661 47075 5695
rect 47501 5661 47535 5695
rect 48237 5661 48271 5695
rect 50445 5661 50479 5695
rect 51273 5661 51307 5695
rect 51917 5661 51951 5695
rect 52745 5661 52779 5695
rect 53389 5661 53423 5695
rect 54125 5661 54159 5695
rect 56333 5661 56367 5695
rect 57989 5661 58023 5695
rect 59553 5661 59587 5695
rect 59737 5661 59771 5695
rect 61485 5661 61519 5695
rect 62957 5661 62991 5695
rect 63141 5661 63175 5695
rect 64889 5661 64923 5695
rect 66361 5661 66395 5695
rect 68293 5661 68327 5695
rect 24133 5593 24167 5627
rect 37013 5593 37047 5627
rect 46305 5593 46339 5627
rect 49617 5593 49651 5627
rect 24685 5525 24719 5559
rect 25145 5525 25179 5559
rect 35725 5525 35759 5559
rect 41705 5525 41739 5559
rect 53297 5525 53331 5559
rect 54769 5525 54803 5559
rect 55873 5525 55907 5559
rect 56149 5525 56183 5559
rect 61301 5525 61335 5559
rect 63325 5525 63359 5559
rect 64705 5525 64739 5559
rect 66545 5525 66579 5559
rect 68109 5525 68143 5559
rect 24409 5185 24443 5219
rect 24869 5185 24903 5219
rect 25605 5185 25639 5219
rect 26065 5185 26099 5219
rect 26433 5185 26467 5219
rect 26525 5185 26559 5219
rect 27261 5185 27295 5219
rect 27721 5185 27755 5219
rect 28273 5185 28307 5219
rect 28457 5185 28491 5219
rect 28897 5183 28931 5217
rect 29561 5185 29595 5219
rect 29653 5185 29687 5219
rect 30113 5185 30147 5219
rect 30665 5185 30699 5219
rect 30849 5185 30883 5219
rect 42993 5185 43027 5219
rect 44189 5185 44223 5219
rect 46305 5185 46339 5219
rect 47225 5185 47259 5219
rect 53113 5185 53147 5219
rect 54769 5185 54803 5219
rect 54953 5185 54987 5219
rect 70225 5185 70259 5219
rect 71697 5185 71731 5219
rect 73445 5185 73479 5219
rect 73537 5185 73571 5219
rect 24225 5117 24259 5151
rect 25421 5117 25455 5151
rect 25881 5117 25915 5151
rect 27077 5117 27111 5151
rect 27537 5117 27571 5151
rect 29101 5117 29135 5151
rect 30297 5117 30331 5151
rect 40417 5117 40451 5151
rect 41061 5117 41095 5151
rect 41521 5117 41555 5151
rect 44557 5117 44591 5151
rect 45385 5117 45419 5151
rect 46121 5117 46155 5151
rect 46581 5117 46615 5151
rect 47501 5117 47535 5151
rect 48145 5117 48179 5151
rect 49157 5117 49191 5151
rect 49801 5117 49835 5151
rect 53297 5117 53331 5151
rect 70409 5117 70443 5151
rect 71881 5117 71915 5151
rect 24685 5049 24719 5083
rect 25789 5049 25823 5083
rect 24593 4981 24627 5015
rect 26249 4981 26283 5015
rect 26709 4981 26743 5015
rect 27445 4981 27479 5015
rect 27905 4981 27939 5015
rect 28089 4981 28123 5015
rect 28733 4981 28767 5015
rect 29377 4981 29411 5015
rect 29929 4981 29963 5015
rect 30481 4981 30515 5015
rect 42165 4981 42199 5015
rect 45109 4981 45143 5015
rect 46029 4981 46063 5015
rect 46489 4981 46523 5015
rect 52929 4981 52963 5015
rect 54585 4981 54619 5015
rect 70041 4981 70075 5015
rect 71513 4981 71547 5015
rect 73261 4981 73295 5015
rect 42625 4777 42659 4811
rect 34161 4641 34195 4675
rect 44097 4641 44131 4675
rect 33977 4573 34011 4607
rect 41245 4573 41279 4607
rect 41981 4573 42015 4607
rect 43361 4573 43395 4607
rect 44281 4573 44315 4607
rect 46673 4573 46707 4607
rect 46843 4575 46877 4609
rect 61209 4573 61243 4607
rect 41889 4437 41923 4471
rect 44005 4437 44039 4471
rect 44465 4437 44499 4471
rect 47041 4437 47075 4471
rect 61117 4437 61151 4471
rect 19717 4097 19751 4131
rect 27629 4097 27663 4131
rect 30849 4097 30883 4131
rect 31309 4097 31343 4131
rect 34713 4097 34747 4131
rect 34897 4097 34931 4131
rect 19533 4029 19567 4063
rect 27905 4029 27939 4063
rect 29745 4029 29779 4063
rect 30389 3893 30423 3927
rect 20269 3689 20303 3723
rect 26065 3689 26099 3723
rect 26249 3689 26283 3723
rect 33057 3689 33091 3723
rect 31861 3621 31895 3655
rect 19441 3553 19475 3587
rect 19993 3553 20027 3587
rect 19165 3485 19199 3519
rect 20177 3485 20211 3519
rect 20821 3485 20855 3519
rect 22569 3485 22603 3519
rect 23489 3485 23523 3519
rect 23581 3485 23615 3519
rect 24961 3485 24995 3519
rect 25237 3485 25271 3519
rect 25513 3485 25547 3519
rect 25789 3485 25823 3519
rect 28089 3485 28123 3519
rect 31217 3485 31251 3519
rect 31677 3485 31711 3519
rect 32229 3485 32263 3519
rect 32873 3485 32907 3519
rect 25881 3417 25915 3451
rect 27721 3417 27755 3451
rect 23213 3349 23247 3383
rect 23305 3349 23339 3383
rect 26086 3349 26120 3383
rect 27629 3349 27663 3383
rect 27905 3349 27939 3383
rect 31401 3349 31435 3383
rect 32413 3349 32447 3383
rect 20545 3145 20579 3179
rect 21281 3145 21315 3179
rect 25881 3145 25915 3179
rect 28089 3145 28123 3179
rect 29469 3145 29503 3179
rect 30205 3145 30239 3179
rect 33517 3145 33551 3179
rect 35081 3145 35115 3179
rect 37013 3145 37047 3179
rect 17877 3077 17911 3111
rect 21122 3077 21156 3111
rect 54585 3077 54619 3111
rect 18153 3009 18187 3043
rect 20637 3009 20671 3043
rect 21373 3009 21407 3043
rect 23121 3009 23155 3043
rect 26157 3009 26191 3043
rect 26709 3009 26743 3043
rect 26893 3009 26927 3043
rect 28549 3009 28583 3043
rect 29101 3009 29135 3043
rect 29561 3009 29595 3043
rect 29745 3009 29779 3043
rect 30021 3009 30055 3043
rect 31585 3009 31619 3043
rect 32045 3009 32079 3043
rect 32965 3009 32999 3043
rect 33333 3009 33367 3043
rect 34069 3009 34103 3043
rect 34529 3009 34563 3043
rect 34897 3009 34931 3043
rect 35909 3009 35943 3043
rect 36277 3009 36311 3043
rect 36829 3009 36863 3043
rect 45937 3009 45971 3043
rect 47501 3009 47535 3043
rect 49065 3009 49099 3043
rect 52929 3009 52963 3043
rect 54217 3009 54251 3043
rect 54677 3009 54711 3043
rect 56241 3009 56275 3043
rect 57805 3009 57839 3043
rect 59461 3009 59495 3043
rect 61209 3009 61243 3043
rect 63233 3009 63267 3043
rect 64797 3009 64831 3043
rect 66453 3009 66487 3043
rect 68109 3009 68143 3043
rect 69857 3009 69891 3043
rect 71421 3009 71455 3043
rect 72893 3009 72927 3043
rect 18981 2941 19015 2975
rect 19165 2941 19199 2975
rect 19901 2941 19935 2975
rect 20913 2941 20947 2975
rect 21005 2941 21039 2975
rect 21741 2941 21775 2975
rect 23765 2941 23799 2975
rect 24317 2941 24351 2975
rect 25329 2941 25363 2975
rect 27077 2941 27111 2975
rect 27537 2941 27571 2975
rect 28917 2941 28951 2975
rect 30297 2941 30331 2975
rect 32229 2941 32263 2975
rect 33885 2941 33919 2975
rect 35817 2941 35851 2975
rect 22477 2873 22511 2907
rect 29929 2873 29963 2907
rect 47685 2873 47719 2907
rect 18429 2805 18463 2839
rect 19809 2805 19843 2839
rect 21465 2805 21499 2839
rect 22385 2805 22419 2839
rect 23213 2805 23247 2839
rect 24961 2805 24995 2839
rect 25973 2805 26007 2839
rect 26525 2805 26559 2839
rect 28365 2805 28399 2839
rect 30941 2805 30975 2839
rect 31493 2805 31527 2839
rect 32873 2805 32907 2839
rect 34253 2805 34287 2839
rect 35173 2805 35207 2839
rect 46121 2805 46155 2839
rect 49249 2805 49283 2839
rect 53113 2805 53147 2839
rect 54861 2805 54895 2839
rect 56425 2805 56459 2839
rect 57989 2805 58023 2839
rect 59645 2805 59679 2839
rect 61393 2805 61427 2839
rect 63049 2805 63083 2839
rect 64613 2805 64647 2839
rect 66269 2805 66303 2839
rect 68293 2805 68327 2839
rect 69673 2805 69707 2839
rect 71237 2805 71271 2839
rect 73077 2805 73111 2839
rect 18245 2601 18279 2635
rect 18981 2601 19015 2635
rect 19901 2601 19935 2635
rect 19993 2601 20027 2635
rect 21373 2601 21407 2635
rect 24133 2601 24167 2635
rect 25237 2601 25271 2635
rect 25329 2601 25363 2635
rect 27537 2601 27571 2635
rect 29285 2601 29319 2635
rect 31677 2533 31711 2567
rect 33149 2533 33183 2567
rect 34253 2533 34287 2567
rect 44373 2533 44407 2567
rect 47041 2533 47075 2567
rect 53941 2533 53975 2567
rect 63233 2533 63267 2567
rect 18429 2465 18463 2499
rect 20637 2465 20671 2499
rect 30941 2465 30975 2499
rect 34989 2465 35023 2499
rect 36553 2465 36587 2499
rect 39221 2465 39255 2499
rect 55597 2465 55631 2499
rect 60749 2465 60783 2499
rect 67465 2465 67499 2499
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 17601 2397 17635 2431
rect 19349 2397 19383 2431
rect 20729 2397 20763 2431
rect 21649 2397 21683 2431
rect 22845 2397 22879 2431
rect 22937 2397 22971 2431
rect 23581 2397 23615 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 26065 2397 26099 2431
rect 26801 2397 26835 2431
rect 27353 2397 27387 2431
rect 28089 2397 28123 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 30021 2397 30055 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 32505 2397 32539 2431
rect 33609 2397 33643 2431
rect 35173 2397 35207 2431
rect 35265 2397 35299 2431
rect 35909 2397 35943 2431
rect 36001 2397 36035 2431
rect 42441 2397 42475 2431
rect 43729 2397 43763 2431
rect 44741 2397 44775 2431
rect 44925 2397 44959 2431
rect 45569 2397 45603 2431
rect 46213 2397 46247 2431
rect 47409 2397 47443 2431
rect 49065 2397 49099 2431
rect 53389 2397 53423 2431
rect 54125 2397 54159 2431
rect 57345 2397 57379 2431
rect 62313 2397 62347 2431
rect 65625 2397 65659 2431
rect 67741 2397 67775 2431
rect 69949 2397 69983 2431
rect 70685 2397 70719 2431
rect 23213 2329 23247 2363
rect 39497 2329 39531 2363
rect 43085 2329 43119 2363
rect 47225 2329 47259 2363
rect 55321 2329 55355 2363
rect 56149 2329 56183 2363
rect 61025 2329 61059 2363
rect 63417 2329 63451 2363
rect 17233 2261 17267 2295
rect 17325 2261 17359 2295
rect 26709 2261 26743 2295
rect 28549 2261 28583 2295
rect 29469 2261 29503 2295
rect 30297 2261 30331 2295
rect 31769 2261 31803 2295
rect 44557 2261 44591 2295
rect 46765 2261 46799 2295
rect 48053 2261 48087 2295
rect 49709 2261 49743 2295
rect 54769 2261 54803 2295
rect 56057 2261 56091 2295
rect 57989 2261 58023 2295
rect 62957 2261 62991 2295
rect 66269 2261 66303 2295
rect 69305 2261 69339 2295
rect 71329 2261 71363 2295
rect 16405 2057 16439 2091
rect 17417 2057 17451 2091
rect 18153 2057 18187 2091
rect 24133 2057 24167 2091
rect 31861 2057 31895 2091
rect 32505 2057 32539 2091
rect 34621 2057 34655 2091
rect 36829 2057 36863 2091
rect 39129 2057 39163 2091
rect 47133 2057 47167 2091
rect 52285 2057 52319 2091
rect 55045 2057 55079 2091
rect 58909 2057 58943 2091
rect 63601 2057 63635 2091
rect 67281 2057 67315 2091
rect 28089 1989 28123 2023
rect 67005 1989 67039 2023
rect 69121 1989 69155 2023
rect 71973 1989 72007 2023
rect 16221 1921 16255 1955
rect 17601 1921 17635 1955
rect 19993 1921 20027 1955
rect 20269 1921 20303 1955
rect 21465 1921 21499 1955
rect 22201 1921 22235 1955
rect 24409 1921 24443 1955
rect 25881 1921 25915 1955
rect 26157 1921 26191 1955
rect 26893 1921 26927 1955
rect 28917 1921 28951 1955
rect 29101 1921 29135 1955
rect 29653 1921 29687 1955
rect 29745 1921 29779 1955
rect 31309 1921 31343 1955
rect 33333 1921 33367 1955
rect 34805 1921 34839 1955
rect 38117 1921 38151 1955
rect 38301 1921 38335 1955
rect 40417 1921 40451 1955
rect 41705 1921 41739 1955
rect 41797 1921 41831 1955
rect 42717 1921 42751 1955
rect 42993 1921 43027 1955
rect 44741 1921 44775 1955
rect 45385 1921 45419 1955
rect 46765 1921 46799 1955
rect 46949 1921 46983 1955
rect 47961 1921 47995 1955
rect 49525 1921 49559 1955
rect 50077 1921 50111 1955
rect 50261 1921 50295 1955
rect 51825 1921 51859 1955
rect 52009 1921 52043 1955
rect 53113 1921 53147 1955
rect 54493 1921 54527 1955
rect 56425 1921 56459 1955
rect 57897 1921 57931 1955
rect 58449 1921 58483 1955
rect 58633 1921 58667 1955
rect 59829 1921 59863 1955
rect 60013 1921 60047 1955
rect 61393 1921 61427 1955
rect 62957 1921 62991 1955
rect 64613 1921 64647 1955
rect 66085 1921 66119 1955
rect 66637 1921 66671 1955
rect 66729 1921 66763 1955
rect 68661 1921 68695 1955
rect 69397 1921 69431 1955
rect 69673 1921 69707 1955
rect 71053 1921 71087 1955
rect 71605 1921 71639 1955
rect 71697 1921 71731 1955
rect 16865 1853 16899 1887
rect 19717 1853 19751 1887
rect 22845 1853 22879 1887
rect 23581 1853 23615 1887
rect 25421 1853 25455 1887
rect 28733 1853 28767 1887
rect 30389 1853 30423 1887
rect 33149 1853 33183 1887
rect 33885 1853 33919 1887
rect 33977 1853 34011 1887
rect 35173 1853 35207 1887
rect 36185 1853 36219 1887
rect 37565 1853 37599 1887
rect 39773 1853 39807 1887
rect 39865 1853 39899 1887
rect 41153 1853 41187 1887
rect 43453 1853 43487 1887
rect 44925 1853 44959 1887
rect 45477 1853 45511 1887
rect 46029 1853 46063 1887
rect 46213 1853 46247 1887
rect 48421 1853 48455 1887
rect 51273 1853 51307 1887
rect 53389 1853 53423 1887
rect 55597 1853 55631 1887
rect 56701 1853 56735 1887
rect 59277 1853 59311 1887
rect 60565 1853 60599 1887
rect 61669 1853 61703 1887
rect 63877 1853 63911 1887
rect 64981 1853 65015 1887
rect 67925 1853 67959 1887
rect 68109 1853 68143 1887
rect 69949 1853 69983 1887
rect 72341 1853 72375 1887
rect 72985 1853 73019 1887
rect 73813 1853 73847 1887
rect 25697 1785 25731 1819
rect 38577 1785 38611 1819
rect 50537 1785 50571 1819
rect 60289 1785 60323 1819
rect 18245 1717 18279 1751
rect 26709 1717 26743 1751
rect 41981 1717 42015 1751
rect 42533 1717 42567 1751
rect 56149 1717 56183 1751
rect 61117 1717 61151 1751
rect 64429 1717 64463 1751
rect 73261 1717 73295 1751
rect 22661 1513 22695 1547
rect 25237 1513 25271 1547
rect 27813 1513 27847 1547
rect 30389 1513 30423 1547
rect 37933 1513 37967 1547
rect 41245 1513 41279 1547
rect 46397 1513 46431 1547
rect 48973 1513 49007 1547
rect 51549 1513 51583 1547
rect 61853 1513 61887 1547
rect 64429 1513 64463 1547
rect 70225 1513 70259 1547
rect 47133 1445 47167 1479
rect 21005 1377 21039 1411
rect 28365 1377 28399 1411
rect 38485 1377 38519 1411
rect 42809 1377 42843 1411
rect 45385 1377 45419 1411
rect 47961 1377 47995 1411
rect 50537 1377 50571 1411
rect 60841 1377 60875 1411
rect 63417 1377 63451 1411
rect 68569 1377 68603 1411
rect 71605 1377 71639 1411
rect 5089 1309 5123 1343
rect 15393 1309 15427 1343
rect 15761 1309 15795 1343
rect 17785 1309 17819 1343
rect 18061 1309 18095 1343
rect 18337 1309 18371 1343
rect 19717 1309 19751 1343
rect 19809 1309 19843 1343
rect 22017 1309 22051 1343
rect 24133 1309 24167 1343
rect 24685 1309 24719 1343
rect 26709 1309 26743 1343
rect 27261 1309 27295 1343
rect 27905 1309 27939 1343
rect 29469 1309 29503 1343
rect 29837 1309 29871 1343
rect 30481 1309 30515 1343
rect 32413 1309 32447 1343
rect 33241 1309 33275 1343
rect 34989 1309 35023 1343
rect 35633 1309 35667 1343
rect 37381 1309 37415 1343
rect 38025 1309 38059 1343
rect 39773 1309 39807 1343
rect 41797 1309 41831 1343
rect 42441 1309 42475 1343
rect 43821 1309 43855 1343
rect 44373 1309 44407 1343
rect 44557 1309 44591 1343
rect 44925 1309 44959 1343
rect 46949 1309 46983 1343
rect 47317 1309 47351 1343
rect 47501 1309 47535 1343
rect 49525 1309 49559 1343
rect 50077 1309 50111 1343
rect 52101 1309 52135 1343
rect 52653 1309 52687 1343
rect 54125 1309 54159 1343
rect 54677 1309 54711 1343
rect 55229 1309 55263 1343
rect 56701 1309 56735 1343
rect 57253 1309 57287 1343
rect 57989 1309 58023 1343
rect 59369 1309 59403 1343
rect 59921 1309 59955 1343
rect 60381 1309 60415 1343
rect 62405 1309 62439 1343
rect 63049 1309 63083 1343
rect 64981 1309 65015 1343
rect 65533 1309 65567 1343
rect 66269 1309 66303 1343
rect 68293 1309 68327 1343
rect 69581 1309 69615 1343
rect 71237 1309 71271 1343
rect 73077 1309 73111 1343
rect 73261 1309 73295 1343
rect 3893 1241 3927 1275
rect 16773 1241 16807 1275
rect 19441 1241 19475 1275
rect 23213 1241 23247 1275
rect 25789 1241 25823 1275
rect 31401 1241 31435 1275
rect 33977 1241 34011 1275
rect 35541 1241 35575 1275
rect 36553 1241 36587 1275
rect 40693 1241 40727 1275
rect 53573 1241 53607 1275
rect 56149 1241 56183 1275
rect 58817 1241 58851 1275
rect 65809 1241 65843 1275
rect 67097 1241 67131 1275
rect 72801 1241 72835 1275
rect 74181 1241 74215 1275
rect 15577 1173 15611 1207
rect 16405 1173 16439 1207
rect 29653 1173 29687 1207
rect 32965 1173 32999 1207
rect 44741 1173 44775 1207
<< metal1 >>
rect 65320 85978 74980 86000
rect 65320 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74980 85978
rect 65320 85904 74980 85926
rect 65320 85434 74980 85456
rect 65320 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 74980 85434
rect 65320 85360 74980 85382
rect 65320 84890 74980 84912
rect 65320 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74980 84890
rect 65320 84816 74980 84838
rect 65320 84346 74980 84368
rect 65320 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 74980 84346
rect 65320 84272 74980 84294
rect 64874 84232 64880 84244
rect 63236 84204 64880 84232
rect 64874 84192 64880 84204
rect 64932 84192 64938 84244
rect 65320 83802 74980 83824
rect 65320 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74980 83802
rect 65320 83728 74980 83750
rect 65320 83258 74980 83280
rect 63236 83144 63264 83256
rect 65320 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 74980 83258
rect 65320 83184 74980 83206
rect 66990 83144 66996 83156
rect 63236 83116 66996 83144
rect 66990 83104 66996 83116
rect 67048 83104 67054 83156
rect 69658 83008 69664 83020
rect 63236 82980 69664 83008
rect 69658 82968 69664 82980
rect 69716 82968 69722 83020
rect 65320 82714 74980 82736
rect 65320 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74980 82714
rect 65320 82640 74980 82662
rect 65320 82170 74980 82192
rect 65320 82118 71858 82170
rect 71910 82118 71922 82170
rect 71974 82118 71986 82170
rect 72038 82118 72050 82170
rect 72102 82118 72114 82170
rect 72166 82118 74980 82170
rect 65320 82096 74980 82118
rect 63236 81784 63264 82052
rect 64874 81784 64880 81796
rect 63236 81756 64880 81784
rect 64874 81744 64880 81756
rect 64932 81744 64938 81796
rect 65320 81626 74980 81648
rect 65320 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74980 81626
rect 65320 81552 74980 81574
rect 65320 81082 74980 81104
rect 63236 80968 63264 81076
rect 65320 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 74980 81082
rect 65320 81008 74980 81030
rect 67082 80968 67088 80980
rect 63236 80940 67088 80968
rect 67082 80928 67088 80940
rect 67140 80928 67146 80980
rect 69750 80832 69756 80844
rect 63236 80804 69756 80832
rect 69750 80792 69756 80804
rect 69808 80792 69814 80844
rect 65320 80538 74980 80560
rect 65320 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74980 80538
rect 65320 80464 74980 80486
rect 65320 79994 74980 80016
rect 65320 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 74980 79994
rect 65320 79920 74980 79942
rect 64874 79880 64880 79892
rect 63236 79852 64880 79880
rect 64874 79840 64880 79852
rect 64932 79840 64938 79892
rect 65320 79450 74980 79472
rect 65320 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74980 79450
rect 65320 79376 74980 79398
rect 65320 78906 74980 78928
rect 63236 78724 63264 78896
rect 65320 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 74980 78906
rect 65320 78832 74980 78854
rect 66438 78724 66444 78736
rect 63236 78696 66444 78724
rect 66438 78684 66444 78696
rect 66496 78684 66502 78736
rect 69934 78656 69940 78668
rect 63236 78628 69940 78656
rect 69934 78616 69940 78628
rect 69992 78616 69998 78668
rect 65320 78362 74980 78384
rect 65320 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74980 78362
rect 65320 78288 74980 78310
rect 65320 77818 74980 77840
rect 65320 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 74980 77818
rect 65320 77744 74980 77766
rect 64874 77704 64880 77716
rect 63236 77676 64880 77704
rect 64874 77664 64880 77676
rect 64932 77664 64938 77716
rect 65320 77274 74980 77296
rect 65320 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74980 77274
rect 65320 77200 74980 77222
rect 65320 76730 74980 76752
rect 63236 76548 63264 76716
rect 65320 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 74980 76730
rect 65320 76656 74980 76678
rect 66254 76548 66260 76560
rect 63236 76520 66260 76548
rect 66254 76508 66260 76520
rect 66312 76508 66318 76560
rect 68462 76480 68468 76492
rect 63236 76452 68468 76480
rect 68462 76440 68468 76452
rect 68520 76440 68526 76492
rect 65320 76186 74980 76208
rect 65320 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74980 76186
rect 65320 76112 74980 76134
rect 65320 75642 74980 75664
rect 65320 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 74980 75642
rect 65320 75568 74980 75590
rect 63236 75188 63264 75512
rect 64874 75188 64880 75200
rect 63236 75160 64880 75188
rect 64874 75148 64880 75160
rect 64932 75148 64938 75200
rect 65320 75098 74980 75120
rect 65320 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74980 75098
rect 65320 75024 74980 75046
rect 67634 74644 67640 74656
rect 63236 74616 67640 74644
rect 63236 74536 63264 74616
rect 67634 74604 67640 74616
rect 67692 74604 67698 74656
rect 65320 74554 74980 74576
rect 65320 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 74980 74554
rect 65320 74480 74980 74502
rect 63236 74100 63264 74284
rect 66162 74100 66168 74112
rect 63236 74072 66168 74100
rect 66162 74060 66168 74072
rect 66220 74060 66226 74112
rect 65320 74010 74980 74032
rect 65320 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74980 74010
rect 65320 73936 74980 73958
rect 65320 73466 74980 73488
rect 65320 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 74980 73466
rect 65320 73392 74980 73414
rect 63236 73216 63264 73332
rect 64874 73216 64880 73228
rect 63236 73188 64880 73216
rect 64874 73176 64880 73188
rect 64932 73176 64938 73228
rect 65320 72922 74980 72944
rect 65320 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74980 72922
rect 65320 72848 74980 72870
rect 65320 72378 74980 72400
rect 63236 72196 63264 72356
rect 65320 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 74980 72378
rect 65320 72304 74980 72326
rect 66346 72196 66352 72208
rect 63236 72168 66352 72196
rect 66346 72156 66352 72168
rect 66404 72156 66410 72208
rect 63236 71924 63264 72104
rect 65978 71924 65984 71936
rect 63236 71896 65984 71924
rect 65978 71884 65984 71896
rect 66036 71884 66042 71936
rect 65320 71834 74980 71856
rect 65320 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74980 71834
rect 65320 71760 74980 71782
rect 65320 71290 74980 71312
rect 65320 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 74980 71290
rect 65320 71216 74980 71238
rect 63236 71148 63816 71176
rect 63788 71108 63816 71148
rect 64874 71108 64880 71120
rect 63788 71080 64880 71108
rect 64874 71068 64880 71080
rect 64932 71068 64938 71120
rect 65320 70746 74980 70768
rect 65320 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74980 70746
rect 65320 70672 74980 70694
rect 65320 70202 74980 70224
rect 63236 70020 63264 70176
rect 65320 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 74980 70202
rect 65320 70128 74980 70150
rect 65518 70020 65524 70032
rect 63236 69992 65524 70020
rect 65518 69980 65524 69992
rect 65576 69980 65582 70032
rect 63236 69612 63264 69924
rect 65320 69658 74980 69680
rect 63678 69612 63684 69624
rect 63236 69584 63684 69612
rect 63678 69572 63684 69584
rect 63736 69572 63742 69624
rect 65320 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74980 69658
rect 65320 69584 74980 69606
rect 65320 69114 74980 69136
rect 65320 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 74980 69114
rect 65320 69040 74980 69062
rect 64874 69000 64880 69012
rect 63144 68972 64880 69000
rect 64874 68960 64880 68972
rect 64932 69000 64938 69012
rect 66530 69000 66536 69012
rect 64932 68972 66536 69000
rect 64932 68960 64938 68972
rect 66530 68960 66536 68972
rect 66588 68960 66594 69012
rect 65320 68570 74980 68592
rect 65320 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74980 68570
rect 65320 68496 74980 68518
rect 65320 68026 74980 68048
rect 63236 67844 63264 67996
rect 65320 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 74980 68026
rect 65320 67952 74980 67974
rect 65886 67844 65892 67856
rect 63236 67816 65892 67844
rect 65886 67804 65892 67816
rect 65944 67804 65950 67856
rect 63236 67640 63264 67744
rect 64598 67640 64604 67652
rect 63236 67612 64604 67640
rect 64598 67600 64604 67612
rect 64656 67600 64662 67652
rect 65320 67482 74980 67504
rect 65320 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74980 67482
rect 65320 67408 74980 67430
rect 65320 66938 74980 66960
rect 65320 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 74980 66938
rect 65320 66864 74980 66886
rect 63236 66484 63264 66792
rect 64874 66484 64880 66496
rect 63236 66456 64880 66484
rect 64874 66444 64880 66456
rect 64932 66444 64938 66496
rect 65320 66394 74980 66416
rect 65320 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74980 66394
rect 65320 66320 74980 66342
rect 65320 65850 74980 65872
rect 63236 65668 63264 65816
rect 65320 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 74980 65850
rect 65320 65776 74980 65798
rect 65426 65668 65432 65680
rect 63236 65640 65432 65668
rect 65426 65628 65432 65640
rect 65484 65628 65490 65680
rect 63236 65396 63264 65564
rect 65702 65396 65708 65408
rect 63236 65368 65708 65396
rect 65702 65356 65708 65368
rect 65760 65356 65766 65408
rect 65320 65306 74980 65328
rect 65320 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74980 65306
rect 65320 65232 74980 65254
rect 65320 64762 74980 64784
rect 65320 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 74980 64762
rect 65320 64688 74980 64710
rect 63236 64308 63264 64612
rect 64874 64308 64880 64320
rect 63236 64280 64880 64308
rect 64874 64268 64880 64280
rect 64932 64268 64938 64320
rect 65320 64218 74980 64240
rect 65320 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74980 64218
rect 65320 64144 74980 64166
rect 65320 63674 74980 63696
rect 63236 63560 63264 63636
rect 65320 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 74980 63674
rect 65320 63600 74980 63622
rect 65334 63560 65340 63572
rect 63236 63532 65340 63560
rect 65334 63520 65340 63532
rect 65392 63520 65398 63572
rect 69014 63424 69020 63436
rect 63236 63396 69020 63424
rect 63236 63384 63264 63396
rect 69014 63384 69020 63396
rect 69072 63384 69078 63436
rect 65320 63130 74980 63152
rect 65320 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74980 63130
rect 65320 63056 74980 63078
rect 65320 62586 74980 62608
rect 65320 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 74980 62586
rect 65320 62512 74980 62534
rect 63236 62132 63264 62432
rect 64874 62132 64880 62144
rect 63236 62104 64880 62132
rect 64874 62092 64880 62104
rect 64932 62092 64938 62144
rect 65320 62042 74980 62064
rect 65320 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74980 62042
rect 65320 61968 74980 61990
rect 65320 61498 74980 61520
rect 63236 61316 63264 61456
rect 65320 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 74980 61498
rect 65320 61424 74980 61446
rect 65242 61316 65248 61328
rect 63236 61288 65248 61316
rect 65242 61276 65248 61288
rect 65300 61276 65306 61328
rect 63236 60908 63264 61204
rect 65320 60954 74980 60976
rect 63586 60908 63592 60920
rect 63236 60880 63592 60908
rect 63586 60868 63592 60880
rect 63644 60868 63650 60920
rect 65320 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74980 60954
rect 65320 60880 74980 60902
rect 65320 60410 74980 60432
rect 65320 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 74980 60410
rect 65320 60336 74980 60358
rect 63144 60268 63816 60296
rect 63144 60252 63172 60268
rect 63788 60228 63816 60268
rect 64874 60228 64880 60240
rect 63788 60200 64880 60228
rect 64874 60188 64880 60200
rect 64932 60188 64938 60240
rect 65320 59866 74980 59888
rect 65320 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74980 59866
rect 65320 59792 74980 59814
rect 65320 59322 74980 59344
rect 63236 59140 63264 59276
rect 65320 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 74980 59322
rect 65320 59248 74980 59270
rect 65150 59140 65156 59152
rect 63236 59112 65156 59140
rect 65150 59100 65156 59112
rect 65208 59100 65214 59152
rect 70762 59072 70768 59084
rect 63236 59044 70768 59072
rect 63236 59024 63264 59044
rect 70762 59032 70768 59044
rect 70820 59032 70826 59084
rect 65320 58778 74980 58800
rect 65320 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74980 58778
rect 65320 58704 74980 58726
rect 65320 58234 74980 58256
rect 65320 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 74980 58234
rect 65320 58160 74980 58182
rect 63236 58052 63264 58072
rect 64874 58052 64880 58064
rect 63236 58024 64880 58052
rect 64874 58012 64880 58024
rect 64932 58012 64938 58064
rect 65320 57690 74980 57712
rect 65320 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74980 57690
rect 65320 57616 74980 57638
rect 65320 57146 74980 57168
rect 63236 57032 63264 57096
rect 65320 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 74980 57146
rect 65320 57072 74980 57094
rect 68094 57032 68100 57044
rect 63236 57004 68100 57032
rect 68094 56992 68100 57004
rect 68152 56992 68158 57044
rect 63236 56692 63264 56844
rect 65794 56692 65800 56704
rect 63236 56664 65800 56692
rect 65794 56652 65800 56664
rect 65852 56652 65858 56704
rect 65320 56602 74980 56624
rect 65320 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74980 56602
rect 65320 56528 74980 56550
rect 65320 56058 74980 56080
rect 65320 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 74980 56058
rect 65320 55984 74980 56006
rect 63236 55604 63264 55892
rect 64874 55604 64880 55616
rect 63236 55576 64880 55604
rect 64874 55564 64880 55576
rect 64932 55564 64938 55616
rect 65320 55514 74980 55536
rect 65320 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74980 55514
rect 65320 55440 74980 55462
rect 65320 54970 74980 54992
rect 65320 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 74980 54970
rect 63236 54788 63264 54916
rect 65320 54896 74980 54918
rect 67542 54788 67548 54800
rect 63236 54760 67548 54788
rect 67542 54748 67548 54760
rect 67600 54748 67606 54800
rect 63144 54652 63172 54664
rect 69106 54652 69112 54664
rect 63144 54624 69112 54652
rect 69106 54612 69112 54624
rect 69164 54612 69170 54664
rect 65320 54426 74980 54448
rect 65320 54374 74210 54426
rect 74262 54374 74274 54426
rect 74326 54374 74338 54426
rect 74390 54374 74402 54426
rect 74454 54374 74466 54426
rect 74518 54374 74980 54426
rect 65320 54352 74980 54374
rect 65320 53882 74980 53904
rect 65320 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 74980 53882
rect 65320 53808 74980 53830
rect 63236 53564 63264 53712
rect 64874 53564 64880 53576
rect 63236 53536 64880 53564
rect 64874 53524 64880 53536
rect 64932 53524 64938 53576
rect 63236 53156 63264 53432
rect 65320 53338 74980 53360
rect 65320 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74980 53338
rect 65320 53264 74980 53286
rect 66898 53156 66904 53168
rect 63236 53128 66904 53156
rect 66898 53116 66904 53128
rect 66956 53116 66962 53168
rect 65320 52794 74980 52816
rect 65320 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 74980 52794
rect 63236 52680 63264 52736
rect 65320 52720 74980 52742
rect 68186 52680 68192 52692
rect 63236 52652 68192 52680
rect 68186 52640 68192 52652
rect 68244 52640 68250 52692
rect 63494 52612 63500 52624
rect 63144 52584 63500 52612
rect 63144 52484 63172 52584
rect 63494 52572 63500 52584
rect 63552 52572 63558 52624
rect 65610 52436 65616 52488
rect 65668 52436 65674 52488
rect 65889 52479 65947 52485
rect 65889 52445 65901 52479
rect 65935 52445 65947 52479
rect 65889 52439 65947 52445
rect 65904 52408 65932 52439
rect 63236 52380 65932 52408
rect 63236 52171 63264 52380
rect 65320 52250 74980 52272
rect 65320 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74980 52250
rect 65320 52176 74980 52198
rect 65610 52136 65616 52148
rect 63604 52108 65616 52136
rect 63250 52080 63632 52108
rect 65610 52096 65616 52108
rect 65668 52096 65674 52148
rect 65320 51706 74980 51728
rect 65320 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 74980 51706
rect 65320 51632 74980 51654
rect 63236 51524 63264 51532
rect 64874 51524 64880 51536
rect 63236 51496 64880 51524
rect 64874 51484 64880 51496
rect 64932 51524 64938 51536
rect 66622 51524 66628 51536
rect 64932 51496 66628 51524
rect 64932 51484 64938 51496
rect 66622 51484 66628 51496
rect 66680 51484 66686 51536
rect 65320 51162 74980 51184
rect 65320 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74980 51162
rect 65320 51088 74980 51110
rect 65320 50618 74980 50640
rect 65320 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 74980 50618
rect 63236 50436 63264 50556
rect 65320 50544 74980 50566
rect 67358 50436 67364 50448
rect 63236 50408 67364 50436
rect 67358 50396 67364 50408
rect 67416 50396 67422 50448
rect 63236 50300 63264 50304
rect 63494 50300 63500 50312
rect 63236 50272 63500 50300
rect 63494 50260 63500 50272
rect 63552 50260 63558 50312
rect 65613 50303 65671 50309
rect 65613 50300 65625 50303
rect 64846 50272 65625 50300
rect 64846 50232 64874 50272
rect 65613 50269 65625 50272
rect 65659 50269 65671 50303
rect 65613 50263 65671 50269
rect 63236 50204 64874 50232
rect 63236 49996 63264 50204
rect 65320 50074 74980 50096
rect 65320 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74980 50074
rect 65320 50000 74980 50022
rect 63250 49643 63632 49671
rect 63604 49620 63632 49643
rect 65613 49623 65671 49629
rect 65613 49620 65625 49623
rect 63604 49592 65625 49620
rect 65613 49589 65625 49592
rect 65659 49589 65671 49623
rect 65613 49583 65671 49589
rect 65320 49530 74980 49552
rect 65320 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 74980 49530
rect 65320 49456 74980 49478
rect 65613 49215 65671 49221
rect 65613 49212 65625 49215
rect 64846 49184 65625 49212
rect 63402 48809 63408 48821
rect 63250 48781 63408 48809
rect 63402 48769 63408 48781
rect 63460 48769 63466 48821
rect 64846 48736 64874 49184
rect 65613 49181 65625 49184
rect 65659 49181 65671 49215
rect 65613 49175 65671 49181
rect 65320 48986 74980 49008
rect 65320 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74980 48986
rect 65320 48912 74980 48934
rect 63604 48729 64874 48736
rect 63250 48708 64874 48729
rect 63250 48701 63632 48708
rect 65320 48442 74980 48464
rect 65320 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 74980 48442
rect 65320 48368 74980 48390
rect 63494 48101 63500 48113
rect 63250 48073 63500 48101
rect 63494 48061 63500 48073
rect 63552 48061 63558 48113
rect 63236 47716 63264 48007
rect 65320 47898 74980 47920
rect 65320 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74980 47898
rect 65320 47824 74980 47846
rect 63862 47716 63868 47728
rect 63236 47688 63868 47716
rect 63862 47676 63868 47688
rect 63920 47676 63926 47728
rect 68554 47512 68560 47524
rect 63144 47484 68560 47512
rect 63144 47379 63172 47484
rect 68554 47472 68560 47484
rect 68612 47472 68618 47524
rect 65320 47354 74980 47376
rect 65320 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 74980 47354
rect 63236 47036 63264 47299
rect 65320 47280 74980 47302
rect 64782 47036 64788 47048
rect 63236 47008 64788 47036
rect 64782 46996 64788 47008
rect 64840 46996 64846 47048
rect 65613 47039 65671 47045
rect 65613 47005 65625 47039
rect 65659 47036 65671 47039
rect 67174 47036 67180 47048
rect 65659 47008 67180 47036
rect 65659 47005 65671 47008
rect 65613 46999 65671 47005
rect 67174 46996 67180 47008
rect 67232 46996 67238 47048
rect 65889 46971 65947 46977
rect 65889 46937 65901 46971
rect 65935 46968 65947 46971
rect 66806 46968 66812 46980
rect 65935 46940 66812 46968
rect 65935 46937 65947 46940
rect 65889 46931 65947 46937
rect 66806 46928 66812 46940
rect 66864 46928 66870 46980
rect 65320 46810 74980 46832
rect 65320 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74980 46810
rect 65320 46736 74980 46758
rect 65320 46266 74980 46288
rect 65320 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 74980 46266
rect 65320 46192 74980 46214
rect 68370 46016 68376 46028
rect 63236 45988 68376 46016
rect 63236 45963 63264 45988
rect 68370 45976 68376 45988
rect 68428 45976 68434 46028
rect 63236 45744 63264 45883
rect 63954 45744 63960 45756
rect 63236 45716 63960 45744
rect 63954 45704 63960 45716
rect 64012 45704 64018 45756
rect 65320 45722 74980 45744
rect 65320 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74980 45722
rect 65320 45648 74980 45670
rect 63250 45268 63632 45269
rect 63862 45268 63868 45280
rect 63250 45241 63868 45268
rect 63604 45240 63868 45241
rect 63862 45228 63868 45240
rect 63920 45228 63926 45280
rect 65320 45178 74980 45200
rect 63236 44860 63264 45175
rect 65320 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 74980 45178
rect 65320 45104 74980 45126
rect 64874 44860 64880 44872
rect 63236 44832 64880 44860
rect 64874 44820 64880 44832
rect 64932 44820 64938 44872
rect 65320 44634 74980 44656
rect 65320 44582 74210 44634
rect 74262 44582 74274 44634
rect 74326 44582 74338 44634
rect 74390 44582 74402 44634
rect 74454 44582 74466 44634
rect 74518 44582 74980 44634
rect 63250 44533 63632 44561
rect 65320 44560 74980 44582
rect 63604 44520 63632 44533
rect 68278 44520 68284 44532
rect 63604 44492 68284 44520
rect 68278 44480 68284 44492
rect 68336 44480 68342 44532
rect 63236 44452 63264 44467
rect 67726 44452 67732 44464
rect 63236 44424 67732 44452
rect 67726 44412 67732 44424
rect 67784 44412 67790 44464
rect 65320 44090 74980 44112
rect 65320 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 74980 44090
rect 65320 44016 74980 44038
rect 64046 43840 64052 43852
rect 63236 43812 64052 43840
rect 64046 43800 64052 43812
rect 64104 43800 64110 43852
rect 65613 43775 65671 43781
rect 65613 43772 65625 43775
rect 63236 43744 65625 43772
rect 63236 43654 63264 43744
rect 65613 43741 65625 43744
rect 65659 43741 65671 43775
rect 65613 43735 65671 43741
rect 65320 43546 74980 43568
rect 65320 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74980 43546
rect 65320 43472 74980 43494
rect 70486 43296 70492 43308
rect 63236 43268 70492 43296
rect 70486 43256 70492 43268
rect 70544 43256 70550 43308
rect 68738 43092 68744 43104
rect 63512 43064 68744 43092
rect 63512 43032 63540 43064
rect 68738 43052 68744 43064
rect 68796 43052 68802 43104
rect 63250 43004 63540 43032
rect 65320 43002 74980 43024
rect 65320 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 74980 43002
rect 65320 42928 74980 42950
rect 66990 42712 66996 42764
rect 67048 42752 67054 42764
rect 68005 42755 68063 42761
rect 68005 42752 68017 42755
rect 67048 42724 68017 42752
rect 67048 42712 67054 42724
rect 68005 42721 68017 42724
rect 68051 42721 68063 42755
rect 68005 42715 68063 42721
rect 65613 42687 65671 42693
rect 65613 42684 65625 42687
rect 63236 42656 65625 42684
rect 63236 42402 63264 42656
rect 65613 42653 65625 42656
rect 65659 42653 65671 42687
rect 65613 42647 65671 42653
rect 68649 42687 68707 42693
rect 68649 42653 68661 42687
rect 68695 42684 68707 42687
rect 70026 42684 70032 42696
rect 68695 42656 70032 42684
rect 68695 42653 68707 42656
rect 68649 42647 68707 42653
rect 70026 42644 70032 42656
rect 70084 42644 70090 42696
rect 65320 42458 74980 42480
rect 65320 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74980 42458
rect 65320 42384 74980 42406
rect 63236 41732 63264 42042
rect 65320 41914 74980 41936
rect 65320 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 74980 41914
rect 65320 41840 74980 41862
rect 67082 41760 67088 41812
rect 67140 41760 67146 41812
rect 65058 41732 65064 41744
rect 63236 41704 65064 41732
rect 65058 41692 65064 41704
rect 65116 41692 65122 41744
rect 67729 41599 67787 41605
rect 67729 41565 67741 41599
rect 67775 41596 67787 41599
rect 70118 41596 70124 41608
rect 67775 41568 70124 41596
rect 67775 41565 67787 41568
rect 67729 41559 67787 41565
rect 70118 41556 70124 41568
rect 70176 41556 70182 41608
rect 65320 41370 74980 41392
rect 65320 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74980 41370
rect 65320 41296 74980 41318
rect 63236 40984 63264 41090
rect 64966 40984 64972 40996
rect 63236 40956 64972 40984
rect 64966 40944 64972 40956
rect 65024 40944 65030 40996
rect 67910 40916 67916 40928
rect 63512 40888 67916 40916
rect 63512 40852 63540 40888
rect 67910 40876 67916 40888
rect 67968 40876 67974 40928
rect 63250 40824 63540 40852
rect 65320 40826 74980 40848
rect 65320 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 74980 40826
rect 65320 40752 74980 40774
rect 66438 40672 66444 40724
rect 66496 40672 66502 40724
rect 67085 40511 67143 40517
rect 67085 40477 67097 40511
rect 67131 40508 67143 40511
rect 69198 40508 69204 40520
rect 67131 40480 69204 40508
rect 67131 40477 67143 40480
rect 67085 40471 67143 40477
rect 69198 40468 69204 40480
rect 69256 40468 69262 40520
rect 65320 40282 74980 40304
rect 65320 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74980 40282
rect 65320 40208 74980 40230
rect 63144 39868 63816 39896
rect 63144 39862 63172 39868
rect 63788 39828 63816 39868
rect 65058 39828 65064 39840
rect 63788 39800 65064 39828
rect 65058 39788 65064 39800
rect 65116 39788 65122 39840
rect 65320 39738 74980 39760
rect 65320 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 74980 39738
rect 65320 39664 74980 39686
rect 65613 39627 65671 39633
rect 65613 39593 65625 39627
rect 65659 39624 65671 39627
rect 66254 39624 66260 39636
rect 65659 39596 66260 39624
rect 65659 39593 65671 39596
rect 65613 39587 65671 39593
rect 66254 39584 66260 39596
rect 66312 39584 66318 39636
rect 66257 39423 66315 39429
rect 66257 39389 66269 39423
rect 66303 39420 66315 39423
rect 67450 39420 67456 39432
rect 66303 39392 67456 39420
rect 66303 39389 66315 39392
rect 66257 39383 66315 39389
rect 67450 39380 67456 39392
rect 67508 39380 67514 39432
rect 65320 39194 74980 39216
rect 65320 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74980 39194
rect 65320 39120 74980 39142
rect 63250 38896 63632 38924
rect 63604 38876 63632 38896
rect 64966 38876 64972 38888
rect 63604 38848 64972 38876
rect 64966 38836 64972 38848
rect 65024 38836 65030 38888
rect 68002 38740 68008 38752
rect 63236 38712 68008 38740
rect 63236 38658 63264 38712
rect 68002 38700 68008 38712
rect 68060 38700 68066 38752
rect 65320 38650 74980 38672
rect 65320 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 74980 38650
rect 65320 38576 74980 38598
rect 65613 38539 65671 38545
rect 65613 38505 65625 38539
rect 65659 38536 65671 38539
rect 67634 38536 67640 38548
rect 65659 38508 67640 38536
rect 65659 38505 65671 38508
rect 65613 38499 65671 38505
rect 67634 38496 67640 38508
rect 67692 38496 67698 38548
rect 66257 38335 66315 38341
rect 66257 38301 66269 38335
rect 66303 38332 66315 38335
rect 66990 38332 66996 38344
rect 66303 38304 66996 38332
rect 66303 38301 66315 38304
rect 66257 38295 66315 38301
rect 66990 38292 66996 38304
rect 67048 38292 67054 38344
rect 65320 38106 74980 38128
rect 65320 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74980 38106
rect 65320 38032 74980 38054
rect 63236 37380 63264 37682
rect 65320 37562 74980 37584
rect 65320 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 74980 37562
rect 65320 37488 74980 37510
rect 65058 37380 65064 37392
rect 63236 37352 65064 37380
rect 65058 37340 65064 37352
rect 65116 37340 65122 37392
rect 66257 37247 66315 37253
rect 66257 37213 66269 37247
rect 66303 37244 66315 37247
rect 67266 37244 67272 37256
rect 66303 37216 67272 37244
rect 66303 37213 66315 37216
rect 66257 37207 66315 37213
rect 67266 37204 67272 37216
rect 67324 37204 67330 37256
rect 65613 37179 65671 37185
rect 65613 37145 65625 37179
rect 65659 37176 65671 37179
rect 66346 37176 66352 37188
rect 65659 37148 66352 37176
rect 65659 37145 65671 37148
rect 65613 37139 65671 37145
rect 66346 37136 66352 37148
rect 66404 37136 66410 37188
rect 65320 37018 74980 37040
rect 65320 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74980 37018
rect 65320 36944 74980 36966
rect 63236 36564 63264 36730
rect 66070 36564 66076 36576
rect 63236 36536 66076 36564
rect 66070 36524 66076 36536
rect 66128 36524 66134 36576
rect 63236 36360 63264 36478
rect 65320 36474 74980 36496
rect 65320 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 74980 36474
rect 65320 36400 74980 36422
rect 63236 36332 64874 36360
rect 64846 36292 64874 36332
rect 65518 36320 65524 36372
rect 65576 36360 65582 36372
rect 65613 36363 65671 36369
rect 65613 36360 65625 36363
rect 65576 36332 65625 36360
rect 65576 36320 65582 36332
rect 65613 36329 65625 36332
rect 65659 36329 65671 36363
rect 65613 36323 65671 36329
rect 69290 36292 69296 36304
rect 64846 36264 69296 36292
rect 69290 36252 69296 36264
rect 69348 36252 69354 36304
rect 66257 36159 66315 36165
rect 66257 36125 66269 36159
rect 66303 36156 66315 36159
rect 66346 36156 66352 36168
rect 66303 36128 66352 36156
rect 66303 36125 66315 36128
rect 66257 36119 66315 36125
rect 66346 36116 66352 36128
rect 66404 36116 66410 36168
rect 65320 35930 74980 35952
rect 65320 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74980 35930
rect 65320 35856 74980 35878
rect 66530 35708 66536 35760
rect 66588 35708 66594 35760
rect 65797 35683 65855 35689
rect 65797 35649 65809 35683
rect 65843 35680 65855 35683
rect 70578 35680 70584 35692
rect 65843 35652 70584 35680
rect 65843 35649 65855 35652
rect 65797 35643 65855 35649
rect 70578 35640 70584 35652
rect 70636 35640 70642 35692
rect 63236 35204 63264 35502
rect 65320 35386 74980 35408
rect 65320 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 74980 35386
rect 65320 35312 74980 35334
rect 65613 35275 65671 35281
rect 65613 35241 65625 35275
rect 65659 35272 65671 35275
rect 65886 35272 65892 35284
rect 65659 35244 65892 35272
rect 65659 35241 65671 35244
rect 65613 35235 65671 35241
rect 65886 35232 65892 35244
rect 65944 35232 65950 35284
rect 64874 35204 64880 35216
rect 63236 35176 64880 35204
rect 64874 35164 64880 35176
rect 64932 35204 64938 35216
rect 65058 35204 65064 35216
rect 64932 35176 65064 35204
rect 64932 35164 64938 35176
rect 65058 35164 65064 35176
rect 65116 35164 65122 35216
rect 66257 35071 66315 35077
rect 66257 35037 66269 35071
rect 66303 35068 66315 35071
rect 67082 35068 67088 35080
rect 66303 35040 67088 35068
rect 66303 35037 66315 35040
rect 66257 35031 66315 35037
rect 67082 35028 67088 35040
rect 67140 35028 67146 35080
rect 65320 34842 74980 34864
rect 65320 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74980 34842
rect 65320 34768 74980 34790
rect 65518 34592 65524 34604
rect 63236 34564 65524 34592
rect 63236 34550 63264 34564
rect 65518 34552 65524 34564
rect 65576 34552 65582 34604
rect 65320 34298 74980 34320
rect 63236 33980 63264 34298
rect 65320 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 74980 34298
rect 65320 34224 74980 34246
rect 66898 34144 66904 34196
rect 66956 34144 66962 34196
rect 64690 33980 64696 33992
rect 63236 33952 64696 33980
rect 64690 33940 64696 33952
rect 64748 33940 64754 33992
rect 65610 33872 65616 33924
rect 65668 33872 65674 33924
rect 65320 33754 74980 33776
rect 65320 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74980 33754
rect 65320 33680 74980 33702
rect 65426 33600 65432 33652
rect 65484 33640 65490 33652
rect 65613 33643 65671 33649
rect 65613 33640 65625 33643
rect 65484 33612 65625 33640
rect 65484 33600 65490 33612
rect 65613 33609 65625 33612
rect 65659 33609 65671 33643
rect 65613 33603 65671 33609
rect 66257 33439 66315 33445
rect 66257 33405 66269 33439
rect 66303 33436 66315 33439
rect 66714 33436 66720 33448
rect 66303 33408 66720 33436
rect 66303 33405 66315 33408
rect 66257 33399 66315 33405
rect 66714 33396 66720 33408
rect 66772 33396 66778 33448
rect 63236 33300 63264 33322
rect 64874 33300 64880 33312
rect 63236 33272 64880 33300
rect 64874 33260 64880 33272
rect 64932 33260 64938 33312
rect 65320 33210 74980 33232
rect 65320 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 74980 33210
rect 65320 33136 74980 33158
rect 65334 33056 65340 33108
rect 65392 33096 65398 33108
rect 65613 33099 65671 33105
rect 65613 33096 65625 33099
rect 65392 33068 65625 33096
rect 65392 33056 65398 33068
rect 65613 33065 65625 33068
rect 65659 33065 65671 33099
rect 65613 33059 65671 33065
rect 66257 32895 66315 32901
rect 66257 32861 66269 32895
rect 66303 32892 66315 32895
rect 66438 32892 66444 32904
rect 66303 32864 66444 32892
rect 66303 32861 66315 32864
rect 66257 32855 66315 32861
rect 66438 32852 66444 32864
rect 66496 32852 66502 32904
rect 65320 32666 74980 32688
rect 65320 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74980 32666
rect 65320 32592 74980 32614
rect 63236 32212 63264 32370
rect 65242 32212 65248 32224
rect 63236 32184 65248 32212
rect 65242 32172 65248 32184
rect 65300 32172 65306 32224
rect 63494 32132 63500 32144
rect 63250 32104 63500 32132
rect 63494 32092 63500 32104
rect 63552 32092 63558 32144
rect 65320 32122 74980 32144
rect 65320 32070 71858 32122
rect 71910 32070 71922 32122
rect 71974 32070 71986 32122
rect 72038 32070 72050 32122
rect 72102 32070 72114 32122
rect 72166 32070 74980 32122
rect 65320 32048 74980 32070
rect 65334 31968 65340 32020
rect 65392 32008 65398 32020
rect 65613 32011 65671 32017
rect 65613 32008 65625 32011
rect 65392 31980 65625 32008
rect 65392 31968 65398 31980
rect 65613 31977 65625 31980
rect 65659 31977 65671 32011
rect 65613 31971 65671 31977
rect 66254 31764 66260 31816
rect 66312 31764 66318 31816
rect 65320 31578 74980 31600
rect 65320 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74980 31578
rect 65320 31504 74980 31526
rect 63236 31124 63264 31142
rect 64874 31124 64880 31136
rect 63236 31096 64880 31124
rect 64874 31084 64880 31096
rect 64932 31084 64938 31136
rect 65320 31034 74980 31056
rect 65320 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 74980 31034
rect 65320 30960 74980 30982
rect 65150 30880 65156 30932
rect 65208 30920 65214 30932
rect 65613 30923 65671 30929
rect 65613 30920 65625 30923
rect 65208 30892 65625 30920
rect 65208 30880 65214 30892
rect 65613 30889 65625 30892
rect 65659 30889 65671 30923
rect 65613 30883 65671 30889
rect 66257 30719 66315 30725
rect 66257 30685 66269 30719
rect 66303 30716 66315 30719
rect 66530 30716 66536 30728
rect 66303 30688 66536 30716
rect 66303 30685 66315 30688
rect 66257 30679 66315 30685
rect 66530 30676 66536 30688
rect 66588 30676 66594 30728
rect 65320 30490 74980 30512
rect 65320 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74980 30490
rect 65320 30416 74980 30438
rect 63236 30036 63264 30190
rect 65334 30036 65340 30048
rect 63236 30008 65340 30036
rect 65334 29996 65340 30008
rect 65392 29996 65398 30048
rect 65320 29946 74980 29968
rect 63236 29628 63264 29938
rect 65320 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 74980 29946
rect 65320 29872 74980 29894
rect 65613 29835 65671 29841
rect 65613 29801 65625 29835
rect 65659 29832 65671 29835
rect 68094 29832 68100 29844
rect 65659 29804 68100 29832
rect 65659 29801 65671 29804
rect 65613 29795 65671 29801
rect 68094 29792 68100 29804
rect 68152 29792 68158 29844
rect 63770 29628 63776 29640
rect 63236 29600 63776 29628
rect 63770 29588 63776 29600
rect 63828 29588 63834 29640
rect 66257 29631 66315 29637
rect 66257 29597 66269 29631
rect 66303 29628 66315 29631
rect 66990 29628 66996 29640
rect 66303 29600 66996 29628
rect 66303 29597 66315 29600
rect 66257 29591 66315 29597
rect 66990 29588 66996 29600
rect 67048 29588 67054 29640
rect 65320 29402 74980 29424
rect 65320 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74980 29402
rect 65320 29328 74980 29350
rect 63236 28676 63264 28962
rect 65320 28858 74980 28880
rect 65320 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 74980 28858
rect 65320 28784 74980 28806
rect 65613 28747 65671 28753
rect 65613 28713 65625 28747
rect 65659 28744 65671 28747
rect 67542 28744 67548 28756
rect 65659 28716 67548 28744
rect 65659 28713 65671 28716
rect 65613 28707 65671 28713
rect 67542 28704 67548 28716
rect 67600 28704 67606 28756
rect 64874 28676 64880 28688
rect 63236 28648 64880 28676
rect 64874 28636 64880 28648
rect 64932 28636 64938 28688
rect 67358 28636 67364 28688
rect 67416 28676 67422 28688
rect 67416 28648 67588 28676
rect 67416 28636 67422 28648
rect 67560 28620 67588 28648
rect 67542 28568 67548 28620
rect 67600 28568 67606 28620
rect 66257 28543 66315 28549
rect 66257 28509 66269 28543
rect 66303 28540 66315 28543
rect 67358 28540 67364 28552
rect 66303 28512 67364 28540
rect 66303 28509 66315 28512
rect 66257 28503 66315 28509
rect 67358 28500 67364 28512
rect 67416 28500 67422 28552
rect 65320 28314 74980 28336
rect 65320 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74980 28314
rect 65320 28240 74980 28262
rect 63236 27860 63264 28010
rect 65886 27860 65892 27872
rect 63236 27832 65892 27860
rect 65886 27820 65892 27832
rect 65944 27820 65950 27872
rect 63494 27772 63500 27784
rect 63250 27744 63500 27772
rect 63494 27732 63500 27744
rect 63552 27732 63558 27784
rect 65320 27770 74980 27792
rect 65320 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 74980 27770
rect 65320 27696 74980 27718
rect 65613 27591 65671 27597
rect 65613 27557 65625 27591
rect 65659 27588 65671 27591
rect 68186 27588 68192 27600
rect 65659 27560 68192 27588
rect 65659 27557 65671 27560
rect 65613 27551 65671 27557
rect 68186 27548 68192 27560
rect 68244 27548 68250 27600
rect 66257 27455 66315 27461
rect 66257 27421 66269 27455
rect 66303 27452 66315 27455
rect 67542 27452 67548 27464
rect 66303 27424 67548 27452
rect 66303 27421 66315 27424
rect 66257 27415 66315 27421
rect 67542 27412 67548 27424
rect 67600 27412 67606 27464
rect 65320 27226 74980 27248
rect 65320 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74980 27226
rect 65320 27152 74980 27174
rect 64874 27112 64880 27124
rect 63236 27084 64880 27112
rect 63236 26782 63264 27084
rect 64874 27072 64880 27084
rect 64932 27112 64938 27124
rect 68094 27112 68100 27124
rect 64932 27084 68100 27112
rect 64932 27072 64938 27084
rect 68094 27072 68100 27084
rect 68152 27072 68158 27124
rect 66622 27004 66628 27056
rect 66680 27004 66686 27056
rect 65797 26979 65855 26985
rect 65797 26945 65809 26979
rect 65843 26976 65855 26979
rect 70670 26976 70676 26988
rect 65843 26948 70676 26976
rect 65843 26945 65855 26948
rect 65797 26939 65855 26945
rect 70670 26936 70676 26948
rect 70728 26936 70734 26988
rect 65320 26682 74980 26704
rect 65320 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 74980 26682
rect 65320 26608 74980 26630
rect 63494 26528 63500 26580
rect 63552 26528 63558 26580
rect 65613 26571 65671 26577
rect 65613 26537 65625 26571
rect 65659 26568 65671 26571
rect 67634 26568 67640 26580
rect 65659 26540 67640 26568
rect 65659 26537 65671 26540
rect 65613 26531 65671 26537
rect 67634 26528 67640 26540
rect 67692 26528 67698 26580
rect 63512 26500 63540 26528
rect 63420 26472 63540 26500
rect 63420 26308 63448 26472
rect 66257 26367 66315 26373
rect 66257 26333 66269 26367
rect 66303 26364 66315 26367
rect 67358 26364 67364 26376
rect 66303 26336 67364 26364
rect 66303 26333 66315 26336
rect 66257 26327 66315 26333
rect 67358 26324 67364 26336
rect 67416 26324 67422 26376
rect 63402 26256 63408 26308
rect 63460 26256 63466 26308
rect 63494 26188 63500 26240
rect 63552 26188 63558 26240
rect 63402 26052 63408 26104
rect 63460 26052 63466 26104
rect 63236 25684 63264 25830
rect 63420 25752 63448 26052
rect 63512 25832 63540 26188
rect 65320 26138 74980 26160
rect 65320 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74980 26138
rect 65320 26064 74980 26086
rect 63586 25984 63592 26036
rect 63644 25984 63650 26036
rect 63604 25832 63632 25984
rect 63494 25780 63500 25832
rect 63552 25780 63558 25832
rect 63586 25780 63592 25832
rect 63644 25780 63650 25832
rect 63678 25752 63684 25764
rect 63420 25724 63684 25752
rect 63678 25712 63684 25724
rect 63736 25712 63742 25764
rect 65426 25684 65432 25696
rect 63236 25656 65432 25684
rect 65426 25644 65432 25656
rect 65484 25644 65490 25696
rect 65320 25594 74980 25616
rect 63236 25480 63264 25578
rect 65320 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 74980 25594
rect 65320 25520 74980 25542
rect 68646 25480 68652 25492
rect 63236 25452 68652 25480
rect 68646 25440 68652 25452
rect 68704 25440 68710 25492
rect 65320 25050 74980 25072
rect 65320 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74980 25050
rect 65320 24976 74980 24998
rect 63236 24324 63264 24602
rect 65320 24506 74980 24528
rect 65320 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 74980 24506
rect 65320 24432 74980 24454
rect 65613 24395 65671 24401
rect 65613 24361 65625 24395
rect 65659 24392 65671 24395
rect 67726 24392 67732 24404
rect 65659 24364 67732 24392
rect 65659 24361 65671 24364
rect 65613 24355 65671 24361
rect 67726 24352 67732 24364
rect 67784 24352 67790 24404
rect 65150 24324 65156 24336
rect 63236 24296 65156 24324
rect 65150 24284 65156 24296
rect 65208 24284 65214 24336
rect 66257 24191 66315 24197
rect 66257 24157 66269 24191
rect 66303 24188 66315 24191
rect 66438 24188 66444 24200
rect 66303 24160 66444 24188
rect 66303 24157 66315 24160
rect 66257 24151 66315 24157
rect 66438 24148 66444 24160
rect 66496 24148 66502 24200
rect 65320 23962 74980 23984
rect 65320 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74980 23962
rect 65320 23888 74980 23910
rect 64966 23808 64972 23860
rect 65024 23848 65030 23860
rect 65613 23851 65671 23857
rect 65613 23848 65625 23851
rect 65024 23820 65625 23848
rect 65024 23808 65030 23820
rect 65613 23817 65625 23820
rect 65659 23817 65671 23851
rect 65613 23811 65671 23817
rect 63236 23508 63264 23650
rect 66257 23647 66315 23653
rect 66257 23613 66269 23647
rect 66303 23644 66315 23647
rect 67634 23644 67640 23656
rect 66303 23616 67640 23644
rect 66303 23613 66315 23616
rect 66257 23607 66315 23613
rect 67634 23604 67640 23616
rect 67692 23604 67698 23656
rect 65518 23508 65524 23520
rect 63236 23480 65524 23508
rect 65518 23468 65524 23480
rect 65576 23468 65582 23520
rect 65320 23418 74980 23440
rect 63236 23304 63264 23398
rect 65320 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 74980 23418
rect 65320 23344 74980 23366
rect 65613 23307 65671 23313
rect 63236 23276 64874 23304
rect 64846 23236 64874 23276
rect 65613 23273 65625 23307
rect 65659 23304 65671 23307
rect 68278 23304 68284 23316
rect 65659 23276 68284 23304
rect 65659 23273 65671 23276
rect 65613 23267 65671 23273
rect 68278 23264 68284 23276
rect 68336 23264 68342 23316
rect 68830 23236 68836 23248
rect 64846 23208 68836 23236
rect 68830 23196 68836 23208
rect 68888 23196 68894 23248
rect 66257 23103 66315 23109
rect 66257 23069 66269 23103
rect 66303 23100 66315 23103
rect 66438 23100 66444 23112
rect 66303 23072 66444 23100
rect 66303 23069 66315 23072
rect 66257 23063 66315 23069
rect 66438 23060 66444 23072
rect 66496 23060 66502 23112
rect 65320 22874 74980 22896
rect 65320 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74980 22874
rect 65320 22800 74980 22822
rect 63236 22148 63264 22422
rect 65320 22330 74980 22352
rect 65320 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 74980 22330
rect 65320 22256 74980 22278
rect 66438 22176 66444 22228
rect 66496 22216 66502 22228
rect 67726 22216 67732 22228
rect 66496 22188 67732 22216
rect 66496 22176 66502 22188
rect 67726 22176 67732 22188
rect 67784 22176 67790 22228
rect 65150 22148 65156 22160
rect 63236 22120 65156 22148
rect 65150 22108 65156 22120
rect 65208 22108 65214 22160
rect 65320 21786 74980 21808
rect 65320 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74980 21786
rect 65320 21712 74980 21734
rect 69382 21536 69388 21548
rect 63604 21508 69388 21536
rect 63604 21484 63632 21508
rect 69382 21496 69388 21508
rect 69440 21496 69446 21548
rect 63250 21456 63632 21484
rect 65320 21242 74980 21264
rect 63236 21128 63264 21218
rect 65320 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 74980 21242
rect 65320 21168 74980 21190
rect 68186 21128 68192 21140
rect 63236 21100 68192 21128
rect 68186 21088 68192 21100
rect 68244 21088 68250 21140
rect 65320 20698 74980 20720
rect 65320 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74980 20698
rect 65320 20624 74980 20646
rect 65150 20244 65156 20256
rect 63236 20216 65156 20244
rect 65150 20204 65156 20216
rect 65208 20204 65214 20256
rect 65320 20154 74980 20176
rect 65320 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 74980 20154
rect 65320 20080 74980 20102
rect 65320 19610 74980 19632
rect 65320 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74980 19610
rect 65320 19536 74980 19558
rect 63236 19156 63264 19290
rect 65058 19156 65064 19168
rect 63236 19128 65064 19156
rect 65058 19116 65064 19128
rect 65116 19116 65122 19168
rect 65320 19066 74980 19088
rect 63236 18952 63264 19038
rect 65320 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 74980 19066
rect 65320 18992 74980 19014
rect 67818 18952 67824 18964
rect 63236 18924 67824 18952
rect 67818 18912 67824 18924
rect 67876 18912 67882 18964
rect 65320 18522 74980 18544
rect 65320 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74980 18522
rect 65320 18448 74980 18470
rect 63236 18000 63264 18062
rect 65150 18000 65156 18012
rect 63236 17972 65156 18000
rect 65150 17960 65156 17972
rect 65208 17960 65214 18012
rect 65320 17978 74980 18000
rect 65320 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 74980 17978
rect 65320 17904 74980 17926
rect 65320 17434 74980 17456
rect 65320 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74980 17434
rect 65320 17360 74980 17382
rect 63236 16980 63264 17110
rect 65610 16980 65616 16992
rect 63236 16952 65616 16980
rect 65610 16940 65616 16952
rect 65668 16940 65674 16992
rect 65320 16890 74980 16912
rect 63236 16640 63264 16858
rect 65320 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 74980 16890
rect 65320 16816 74980 16838
rect 63402 16640 63408 16652
rect 63236 16612 63408 16640
rect 63402 16600 63408 16612
rect 63460 16600 63466 16652
rect 63402 16396 63408 16448
rect 63460 16436 63466 16448
rect 63770 16436 63776 16448
rect 63460 16408 63776 16436
rect 63460 16396 63466 16408
rect 63770 16396 63776 16408
rect 63828 16396 63834 16448
rect 65320 16346 74980 16368
rect 65320 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74980 16346
rect 65320 16272 74980 16294
rect 63236 15620 63264 15882
rect 65320 15802 74980 15824
rect 65320 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 74980 15802
rect 65320 15728 74980 15750
rect 65150 15620 65156 15632
rect 63236 15592 65156 15620
rect 65150 15580 65156 15592
rect 65208 15580 65214 15632
rect 65320 15258 74980 15280
rect 65320 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74980 15258
rect 65320 15184 74980 15206
rect 63236 14804 63264 14930
rect 64966 14804 64972 14816
rect 63236 14776 64972 14804
rect 64966 14764 64972 14776
rect 65024 14764 65030 14816
rect 65320 14714 74980 14736
rect 63236 14600 63264 14678
rect 65320 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 74980 14714
rect 65320 14640 74980 14662
rect 67634 14600 67640 14612
rect 63236 14572 67640 14600
rect 67634 14560 67640 14572
rect 67692 14560 67698 14612
rect 65320 14170 74980 14192
rect 65320 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74980 14170
rect 65320 14096 74980 14118
rect 65150 13716 65156 13728
rect 63250 13688 65156 13716
rect 65150 13676 65156 13688
rect 65208 13676 65214 13728
rect 65320 13626 74980 13648
rect 65320 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 74980 13626
rect 65320 13552 74980 13574
rect 65320 13082 74980 13104
rect 65320 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74980 13082
rect 65320 13008 74980 13030
rect 64874 12764 64880 12776
rect 63250 12736 64880 12764
rect 64874 12724 64880 12736
rect 64932 12724 64938 12776
rect 67726 12628 67732 12640
rect 63236 12600 67732 12628
rect 63236 12498 63264 12600
rect 67726 12588 67732 12600
rect 67784 12588 67790 12640
rect 65320 12538 74980 12560
rect 65320 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 74980 12538
rect 65320 12464 74980 12486
rect 63402 12112 63408 12164
rect 63460 12152 63466 12164
rect 63862 12152 63868 12164
rect 63460 12124 63868 12152
rect 63460 12112 63466 12124
rect 63862 12112 63868 12124
rect 63920 12112 63926 12164
rect 65320 11994 74980 12016
rect 65320 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74980 11994
rect 65320 11920 74980 11942
rect 63494 11840 63500 11892
rect 63552 11880 63558 11892
rect 63770 11880 63776 11892
rect 63552 11852 63776 11880
rect 63552 11840 63558 11852
rect 63770 11840 63776 11852
rect 63828 11840 63834 11892
rect 63236 11268 63264 11522
rect 65320 11450 74980 11472
rect 65320 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 74980 11450
rect 65320 11376 74980 11398
rect 65150 11268 65156 11280
rect 63236 11240 65156 11268
rect 65150 11228 65156 11240
rect 65208 11228 65214 11280
rect 64046 11024 64052 11076
rect 64104 11064 64110 11076
rect 66806 11064 66812 11076
rect 64104 11036 66812 11064
rect 64104 11024 64110 11036
rect 66806 11024 66812 11036
rect 66864 11024 66870 11076
rect 65320 10906 74980 10928
rect 65320 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74980 10906
rect 65320 10832 74980 10854
rect 63236 10452 63264 10570
rect 64874 10452 64880 10464
rect 63236 10424 64880 10452
rect 64874 10412 64880 10424
rect 64932 10412 64938 10464
rect 65320 10362 74980 10384
rect 63402 10332 63408 10344
rect 63250 10304 63408 10332
rect 63402 10292 63408 10304
rect 63460 10292 63466 10344
rect 65320 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 74980 10362
rect 65320 10288 74980 10310
rect 65320 9818 74980 9840
rect 65320 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74980 9818
rect 65320 9744 74980 9766
rect 65150 9364 65156 9376
rect 63236 9336 65156 9364
rect 65150 9324 65156 9336
rect 65208 9324 65214 9376
rect 65320 9274 74980 9296
rect 65320 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 74980 9274
rect 65320 9200 74980 9222
rect 65320 8730 74980 8752
rect 65320 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74980 8730
rect 65320 8656 74980 8678
rect 65320 8186 74980 8208
rect 65320 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 74980 8186
rect 65320 8112 74980 8134
rect 62942 7828 62948 7880
rect 63000 7868 63006 7880
rect 65610 7868 65616 7880
rect 63000 7840 65616 7868
rect 63000 7828 63006 7840
rect 65610 7828 65616 7840
rect 65668 7828 65674 7880
rect 52270 7760 52276 7812
rect 52328 7800 52334 7812
rect 60734 7800 60740 7812
rect 52328 7772 60740 7800
rect 52328 7760 52334 7772
rect 60734 7760 60740 7772
rect 60792 7760 60798 7812
rect 61654 7760 61660 7812
rect 61712 7800 61718 7812
rect 64598 7800 64604 7812
rect 61712 7772 64604 7800
rect 61712 7760 61718 7772
rect 64598 7760 64604 7772
rect 64656 7760 64662 7812
rect 43530 7692 43536 7744
rect 43588 7732 43594 7744
rect 62758 7732 62764 7744
rect 43588 7704 62764 7732
rect 43588 7692 43594 7704
rect 62758 7692 62764 7704
rect 62816 7692 62822 7744
rect 62850 7692 62856 7744
rect 62908 7732 62914 7744
rect 64966 7732 64972 7744
rect 62908 7704 64972 7732
rect 62908 7692 62914 7704
rect 64966 7692 64972 7704
rect 65024 7692 65030 7744
rect 48038 7624 48044 7676
rect 48096 7664 48102 7676
rect 48096 7636 48314 7664
rect 48096 7624 48102 7636
rect 24578 7556 24584 7608
rect 24636 7596 24642 7608
rect 24636 7568 41414 7596
rect 24636 7556 24642 7568
rect 41386 7460 41414 7568
rect 48286 7528 48314 7636
rect 55582 7624 55588 7676
rect 55640 7664 55646 7676
rect 63402 7664 63408 7676
rect 55640 7636 63408 7664
rect 55640 7624 55646 7636
rect 63402 7624 63408 7636
rect 63460 7624 63466 7676
rect 65320 7642 74980 7664
rect 54846 7556 54852 7608
rect 54904 7596 54910 7608
rect 65058 7596 65064 7608
rect 54904 7568 65064 7596
rect 54904 7556 54910 7568
rect 65058 7556 65064 7568
rect 65116 7556 65122 7608
rect 65320 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74980 7642
rect 65320 7568 74980 7590
rect 48286 7500 57974 7528
rect 54662 7460 54668 7472
rect 41386 7432 54668 7460
rect 54662 7420 54668 7432
rect 54720 7420 54726 7472
rect 57946 7392 57974 7500
rect 60734 7488 60740 7540
rect 60792 7528 60798 7540
rect 67818 7528 67824 7540
rect 60792 7500 67824 7528
rect 60792 7488 60798 7500
rect 67818 7488 67824 7500
rect 67876 7488 67882 7540
rect 62758 7420 62764 7472
rect 62816 7460 62822 7472
rect 68094 7460 68100 7472
rect 62816 7432 68100 7460
rect 62816 7420 62822 7432
rect 68094 7420 68100 7432
rect 68152 7420 68158 7472
rect 63494 7392 63500 7404
rect 57946 7364 63500 7392
rect 63494 7352 63500 7364
rect 63552 7352 63558 7404
rect 60734 7284 60740 7336
rect 60792 7324 60798 7336
rect 65702 7324 65708 7336
rect 60792 7296 65708 7324
rect 60792 7284 60798 7296
rect 65702 7284 65708 7296
rect 65760 7284 65766 7336
rect 62666 7216 62672 7268
rect 62724 7256 62730 7268
rect 65794 7256 65800 7268
rect 62724 7228 65800 7256
rect 62724 7216 62730 7228
rect 65794 7216 65800 7228
rect 65852 7216 65858 7268
rect 59078 7148 59084 7200
rect 59136 7188 59142 7200
rect 65886 7188 65892 7200
rect 59136 7160 65892 7188
rect 59136 7148 59142 7160
rect 65886 7148 65892 7160
rect 65944 7148 65950 7200
rect 60458 7080 60464 7132
rect 60516 7120 60522 7132
rect 64598 7120 64604 7132
rect 60516 7092 64604 7120
rect 60516 7080 60522 7092
rect 64598 7080 64604 7092
rect 64656 7080 64662 7132
rect 65320 7098 74980 7120
rect 65058 7052 65064 7064
rect 57946 7024 65064 7052
rect 55766 6944 55772 6996
rect 55824 6984 55830 6996
rect 57946 6984 57974 7024
rect 65058 7012 65064 7024
rect 65116 7012 65122 7064
rect 65320 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 74980 7098
rect 65320 7024 74980 7046
rect 55824 6956 57974 6984
rect 55824 6944 55830 6956
rect 54662 6876 54668 6928
rect 54720 6916 54726 6928
rect 54720 6888 55996 6916
rect 54720 6876 54726 6888
rect 46106 6808 46112 6860
rect 46164 6848 46170 6860
rect 55858 6848 55864 6860
rect 46164 6820 55864 6848
rect 46164 6808 46170 6820
rect 55858 6808 55864 6820
rect 55916 6808 55922 6860
rect 55968 6848 55996 6888
rect 61010 6876 61016 6928
rect 61068 6916 61074 6928
rect 61068 6888 65012 6916
rect 61068 6876 61074 6888
rect 60550 6848 60556 6860
rect 55968 6820 60556 6848
rect 60550 6808 60556 6820
rect 60608 6808 60614 6860
rect 61378 6808 61384 6860
rect 61436 6848 61442 6860
rect 64874 6848 64880 6860
rect 61436 6820 64880 6848
rect 61436 6808 61442 6820
rect 64874 6808 64880 6820
rect 64932 6808 64938 6860
rect 64984 6848 65012 6888
rect 65720 6888 66852 6916
rect 65720 6848 65748 6888
rect 64984 6820 65748 6848
rect 65794 6808 65800 6860
rect 65852 6848 65858 6860
rect 66714 6848 66720 6860
rect 65852 6820 66720 6848
rect 65852 6808 65858 6820
rect 66714 6808 66720 6820
rect 66772 6808 66778 6860
rect 66824 6848 66852 6888
rect 69382 6848 69388 6860
rect 66824 6820 69388 6848
rect 69382 6808 69388 6820
rect 69440 6808 69446 6860
rect 48866 6740 48872 6792
rect 48924 6780 48930 6792
rect 63678 6780 63684 6792
rect 48924 6752 63684 6780
rect 48924 6740 48930 6752
rect 63678 6740 63684 6752
rect 63736 6740 63742 6792
rect 64966 6740 64972 6792
rect 65024 6780 65030 6792
rect 67910 6780 67916 6792
rect 65024 6752 67916 6780
rect 65024 6740 65030 6752
rect 67910 6740 67916 6752
rect 67968 6740 67974 6792
rect 42610 6672 42616 6724
rect 42668 6712 42674 6724
rect 42668 6684 64736 6712
rect 42668 6672 42674 6684
rect 27522 6604 27528 6656
rect 27580 6644 27586 6656
rect 61378 6644 61384 6656
rect 27580 6616 61384 6644
rect 27580 6604 27586 6616
rect 61378 6604 61384 6616
rect 61436 6604 61442 6656
rect 23290 6536 23296 6588
rect 23348 6576 23354 6588
rect 62942 6576 62948 6588
rect 23348 6548 62948 6576
rect 23348 6536 23354 6548
rect 62942 6536 62948 6548
rect 63000 6536 63006 6588
rect 64708 6576 64736 6684
rect 65702 6672 65708 6724
rect 65760 6712 65766 6724
rect 67082 6712 67088 6724
rect 65760 6684 67088 6712
rect 65760 6672 65766 6684
rect 67082 6672 67088 6684
rect 67140 6672 67146 6724
rect 65058 6604 65064 6656
rect 65116 6644 65122 6656
rect 68830 6644 68836 6656
rect 65116 6616 68836 6644
rect 65116 6604 65122 6616
rect 68830 6604 68836 6616
rect 68888 6604 68894 6656
rect 64966 6576 64972 6588
rect 64708 6548 64972 6576
rect 64966 6536 64972 6548
rect 65024 6536 65030 6588
rect 65320 6554 74980 6576
rect 28902 6468 28908 6520
rect 28960 6508 28966 6520
rect 46382 6508 46388 6520
rect 28960 6480 46388 6508
rect 28960 6468 28966 6480
rect 46382 6468 46388 6480
rect 46440 6468 46446 6520
rect 51718 6468 51724 6520
rect 51776 6508 51782 6520
rect 55766 6508 55772 6520
rect 51776 6480 55772 6508
rect 51776 6468 51782 6480
rect 55766 6468 55772 6480
rect 55824 6468 55830 6520
rect 55858 6468 55864 6520
rect 55916 6508 55922 6520
rect 64690 6508 64696 6520
rect 55916 6480 64696 6508
rect 55916 6468 55922 6480
rect 64690 6468 64696 6480
rect 64748 6468 64754 6520
rect 65320 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74980 6554
rect 65320 6480 74980 6502
rect 24762 6400 24768 6452
rect 24820 6440 24826 6452
rect 60826 6440 60832 6452
rect 24820 6412 60832 6440
rect 24820 6400 24826 6412
rect 60826 6400 60832 6412
rect 60884 6400 60890 6452
rect 61010 6400 61016 6452
rect 61068 6440 61074 6452
rect 63402 6440 63408 6452
rect 61068 6412 63408 6440
rect 61068 6400 61074 6412
rect 63402 6400 63408 6412
rect 63460 6400 63466 6452
rect 63678 6400 63684 6452
rect 63736 6440 63742 6452
rect 66254 6440 66260 6452
rect 63736 6412 66260 6440
rect 63736 6400 63742 6412
rect 66254 6400 66260 6412
rect 66312 6400 66318 6452
rect 32950 6332 32956 6384
rect 33008 6372 33014 6384
rect 48222 6372 48228 6384
rect 33008 6344 48228 6372
rect 33008 6332 33014 6344
rect 48222 6332 48228 6344
rect 48280 6332 48286 6384
rect 54846 6332 54852 6384
rect 54904 6372 54910 6384
rect 67726 6372 67732 6384
rect 54904 6344 67732 6372
rect 54904 6332 54910 6344
rect 67726 6332 67732 6344
rect 67784 6332 67790 6384
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 32858 6304 32864 6316
rect 23716 6276 32864 6304
rect 23716 6264 23722 6276
rect 32858 6264 32864 6276
rect 32916 6264 32922 6316
rect 51074 6264 51080 6316
rect 51132 6304 51138 6316
rect 63954 6304 63960 6316
rect 51132 6276 63960 6304
rect 51132 6264 51138 6276
rect 63954 6264 63960 6276
rect 64012 6264 64018 6316
rect 64966 6264 64972 6316
rect 65024 6304 65030 6316
rect 68646 6304 68652 6316
rect 65024 6276 68652 6304
rect 65024 6264 65030 6276
rect 68646 6264 68652 6276
rect 68704 6264 68710 6316
rect 27062 6196 27068 6248
rect 27120 6236 27126 6248
rect 45646 6236 45652 6248
rect 27120 6208 45652 6236
rect 27120 6196 27126 6208
rect 45646 6196 45652 6208
rect 45704 6196 45710 6248
rect 48130 6196 48136 6248
rect 48188 6236 48194 6248
rect 48188 6208 51212 6236
rect 48188 6196 48194 6208
rect 24946 6128 24952 6180
rect 25004 6168 25010 6180
rect 44910 6168 44916 6180
rect 25004 6140 44916 6168
rect 25004 6128 25010 6140
rect 44910 6128 44916 6140
rect 44968 6128 44974 6180
rect 47026 6128 47032 6180
rect 47084 6168 47090 6180
rect 51074 6168 51080 6180
rect 47084 6140 51080 6168
rect 47084 6128 47090 6140
rect 51074 6128 51080 6140
rect 51132 6128 51138 6180
rect 51184 6168 51212 6208
rect 53282 6196 53288 6248
rect 53340 6236 53346 6248
rect 57422 6236 57428 6248
rect 53340 6208 57428 6236
rect 53340 6196 53346 6208
rect 57422 6196 57428 6208
rect 57480 6196 57486 6248
rect 57514 6196 57520 6248
rect 57572 6236 57578 6248
rect 60458 6236 60464 6248
rect 57572 6208 60464 6236
rect 57572 6196 57578 6208
rect 60458 6196 60464 6208
rect 60516 6196 60522 6248
rect 60642 6196 60648 6248
rect 60700 6236 60706 6248
rect 63862 6236 63868 6248
rect 60700 6208 63868 6236
rect 60700 6196 60706 6208
rect 63862 6196 63868 6208
rect 63920 6196 63926 6248
rect 64690 6196 64696 6248
rect 64748 6236 64754 6248
rect 66990 6236 66996 6248
rect 64748 6208 66996 6236
rect 64748 6196 64754 6208
rect 66990 6196 66996 6208
rect 67048 6196 67054 6248
rect 63770 6168 63776 6180
rect 51184 6140 63776 6168
rect 63770 6128 63776 6140
rect 63828 6128 63834 6180
rect 64598 6128 64604 6180
rect 64656 6168 64662 6180
rect 68370 6168 68376 6180
rect 64656 6140 68376 6168
rect 64656 6128 64662 6140
rect 68370 6128 68376 6140
rect 68428 6128 68434 6180
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 34882 6100 34888 6112
rect 26200 6072 34888 6100
rect 26200 6060 26206 6072
rect 34882 6060 34888 6072
rect 34940 6060 34946 6112
rect 45554 6060 45560 6112
rect 45612 6100 45618 6112
rect 55674 6100 55680 6112
rect 45612 6072 55680 6100
rect 45612 6060 45618 6072
rect 55674 6060 55680 6072
rect 55732 6060 55738 6112
rect 55858 6060 55864 6112
rect 55916 6100 55922 6112
rect 62850 6100 62856 6112
rect 55916 6072 62856 6100
rect 55916 6060 55922 6072
rect 62850 6060 62856 6072
rect 62908 6060 62914 6112
rect 63402 6060 63408 6112
rect 63460 6100 63466 6112
rect 68186 6100 68192 6112
rect 63460 6072 68192 6100
rect 63460 6060 63466 6072
rect 68186 6060 68192 6072
rect 68244 6060 68250 6112
rect 1012 6010 74980 6032
rect 1012 5958 1858 6010
rect 1910 5958 1922 6010
rect 1974 5958 1986 6010
rect 2038 5958 2050 6010
rect 2102 5958 2114 6010
rect 2166 5958 11858 6010
rect 11910 5958 11922 6010
rect 11974 5958 11986 6010
rect 12038 5958 12050 6010
rect 12102 5958 12114 6010
rect 12166 5958 21858 6010
rect 21910 5958 21922 6010
rect 21974 5958 21986 6010
rect 22038 5958 22050 6010
rect 22102 5958 22114 6010
rect 22166 5958 31858 6010
rect 31910 5958 31922 6010
rect 31974 5958 31986 6010
rect 32038 5958 32050 6010
rect 32102 5958 32114 6010
rect 32166 5958 41858 6010
rect 41910 5958 41922 6010
rect 41974 5958 41986 6010
rect 42038 5958 42050 6010
rect 42102 5958 42114 6010
rect 42166 5958 51858 6010
rect 51910 5958 51922 6010
rect 51974 5958 51986 6010
rect 52038 5958 52050 6010
rect 52102 5958 52114 6010
rect 52166 5958 61858 6010
rect 61910 5958 61922 6010
rect 61974 5958 61986 6010
rect 62038 5958 62050 6010
rect 62102 5958 62114 6010
rect 62166 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 74980 6010
rect 1012 5936 74980 5958
rect 23658 5856 23664 5908
rect 23716 5856 23722 5908
rect 23768 5868 24900 5896
rect 23290 5720 23296 5772
rect 23348 5720 23354 5772
rect 23768 5769 23796 5868
rect 24872 5828 24900 5868
rect 26142 5856 26148 5908
rect 26200 5856 26206 5908
rect 29546 5856 29552 5908
rect 29604 5896 29610 5908
rect 47486 5896 47492 5908
rect 29604 5868 47492 5896
rect 29604 5856 29610 5868
rect 47486 5856 47492 5868
rect 47544 5856 47550 5908
rect 48130 5856 48136 5908
rect 48188 5856 48194 5908
rect 48866 5856 48872 5908
rect 48924 5856 48930 5908
rect 51077 5899 51135 5905
rect 51077 5865 51089 5899
rect 51123 5896 51135 5899
rect 53282 5896 53288 5908
rect 51123 5868 53288 5896
rect 51123 5865 51135 5868
rect 51077 5859 51135 5865
rect 53282 5856 53288 5868
rect 53340 5856 53346 5908
rect 54021 5899 54079 5905
rect 54021 5865 54033 5899
rect 54067 5896 54079 5899
rect 54067 5868 57376 5896
rect 54067 5865 54079 5868
rect 54021 5859 54079 5865
rect 55858 5828 55864 5840
rect 24872 5800 55864 5828
rect 55858 5788 55864 5800
rect 55916 5788 55922 5840
rect 57348 5828 57376 5868
rect 57422 5856 57428 5908
rect 57480 5896 57486 5908
rect 60826 5896 60832 5908
rect 57480 5868 60832 5896
rect 57480 5856 57486 5868
rect 60826 5856 60832 5868
rect 60884 5856 60890 5908
rect 62574 5896 62580 5908
rect 60936 5868 62580 5896
rect 60936 5828 60964 5868
rect 62574 5856 62580 5868
rect 62632 5856 62638 5908
rect 62758 5856 62764 5908
rect 62816 5896 62822 5908
rect 63402 5896 63408 5908
rect 62816 5868 63408 5896
rect 62816 5856 62822 5868
rect 63402 5856 63408 5868
rect 63460 5856 63466 5908
rect 63770 5856 63776 5908
rect 63828 5896 63834 5908
rect 65242 5896 65248 5908
rect 63828 5868 65248 5896
rect 63828 5856 63834 5868
rect 65242 5856 65248 5868
rect 65300 5856 65306 5908
rect 67634 5828 67640 5840
rect 57348 5800 60964 5828
rect 64156 5800 67640 5828
rect 23753 5763 23811 5769
rect 23753 5729 23765 5763
rect 23799 5729 23811 5763
rect 23753 5723 23811 5729
rect 24305 5763 24363 5769
rect 24305 5729 24317 5763
rect 24351 5760 24363 5763
rect 24578 5760 24584 5772
rect 24351 5732 24584 5760
rect 24351 5729 24363 5732
rect 24305 5723 24363 5729
rect 24578 5720 24584 5732
rect 24636 5720 24642 5772
rect 24762 5720 24768 5772
rect 24820 5720 24826 5772
rect 25038 5720 25044 5772
rect 25096 5760 25102 5772
rect 32214 5760 32220 5772
rect 25096 5732 32220 5760
rect 25096 5720 25102 5732
rect 32214 5720 32220 5732
rect 32272 5720 32278 5772
rect 33870 5720 33876 5772
rect 33928 5760 33934 5772
rect 33928 5732 44864 5760
rect 33928 5720 33934 5732
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 23937 5695 23995 5701
rect 23937 5692 23949 5695
rect 23523 5664 23949 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 23937 5661 23949 5664
rect 23983 5692 23995 5695
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 23983 5664 24501 5692
rect 23983 5661 23995 5664
rect 23937 5655 23995 5661
rect 24489 5661 24501 5664
rect 24535 5692 24547 5695
rect 24949 5695 25007 5701
rect 24949 5692 24961 5695
rect 24535 5664 24961 5692
rect 24535 5661 24547 5664
rect 24489 5655 24547 5661
rect 24949 5661 24961 5664
rect 24995 5692 25007 5695
rect 25590 5692 25596 5704
rect 24995 5664 25596 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 25958 5652 25964 5704
rect 26016 5652 26022 5704
rect 40402 5652 40408 5704
rect 40460 5652 40466 5704
rect 41598 5652 41604 5704
rect 41656 5692 41662 5704
rect 42337 5695 42395 5701
rect 42337 5692 42349 5695
rect 41656 5664 42349 5692
rect 41656 5652 41662 5664
rect 42337 5661 42349 5664
rect 42383 5661 42395 5695
rect 42337 5655 42395 5661
rect 43530 5652 43536 5704
rect 43588 5652 43594 5704
rect 43622 5652 43628 5704
rect 43680 5692 43686 5704
rect 43809 5695 43867 5701
rect 43809 5692 43821 5695
rect 43680 5664 43821 5692
rect 43680 5652 43686 5664
rect 43809 5661 43821 5664
rect 43855 5661 43867 5695
rect 43809 5655 43867 5661
rect 44453 5695 44511 5701
rect 44453 5661 44465 5695
rect 44499 5692 44511 5695
rect 44634 5692 44640 5704
rect 44499 5664 44640 5692
rect 44499 5661 44511 5664
rect 44453 5655 44511 5661
rect 44634 5652 44640 5664
rect 44692 5652 44698 5704
rect 44836 5692 44864 5732
rect 44910 5720 44916 5772
rect 44968 5720 44974 5772
rect 48961 5763 49019 5769
rect 48961 5760 48973 5763
rect 45020 5732 48973 5760
rect 45020 5692 45048 5732
rect 48961 5729 48973 5732
rect 49007 5729 49019 5763
rect 48961 5723 49019 5729
rect 49786 5720 49792 5772
rect 49844 5760 49850 5772
rect 51718 5760 51724 5772
rect 49844 5732 51724 5760
rect 49844 5720 49850 5732
rect 51718 5720 51724 5732
rect 51776 5720 51782 5772
rect 55214 5720 55220 5772
rect 55272 5720 55278 5772
rect 56502 5720 56508 5772
rect 56560 5720 56566 5772
rect 57790 5720 57796 5772
rect 57848 5720 57854 5772
rect 58158 5720 58164 5772
rect 58216 5720 58222 5772
rect 59357 5763 59415 5769
rect 59357 5729 59369 5763
rect 59403 5760 59415 5763
rect 59446 5760 59452 5772
rect 59403 5732 59452 5760
rect 59403 5729 59415 5732
rect 59357 5723 59415 5729
rect 59446 5720 59452 5732
rect 59504 5720 59510 5772
rect 59556 5732 61148 5760
rect 44836 5664 45048 5692
rect 45554 5652 45560 5704
rect 45612 5652 45618 5704
rect 45646 5652 45652 5704
rect 45704 5652 45710 5704
rect 46382 5652 46388 5704
rect 46440 5652 46446 5704
rect 47026 5652 47032 5704
rect 47084 5652 47090 5704
rect 47486 5652 47492 5704
rect 47544 5652 47550 5704
rect 48222 5652 48228 5704
rect 48280 5652 48286 5704
rect 50430 5652 50436 5704
rect 50488 5652 50494 5704
rect 51258 5652 51264 5704
rect 51316 5652 51322 5704
rect 51905 5695 51963 5701
rect 51905 5661 51917 5695
rect 51951 5692 51963 5695
rect 52270 5692 52276 5704
rect 51951 5664 52276 5692
rect 51951 5661 51963 5664
rect 51905 5655 51963 5661
rect 52270 5652 52276 5664
rect 52328 5652 52334 5704
rect 52733 5695 52791 5701
rect 52733 5661 52745 5695
rect 52779 5661 52791 5695
rect 52733 5655 52791 5661
rect 24121 5627 24179 5633
rect 24121 5593 24133 5627
rect 24167 5624 24179 5627
rect 24167 5596 31754 5624
rect 24167 5593 24179 5596
rect 24121 5587 24179 5593
rect 24673 5559 24731 5565
rect 24673 5525 24685 5559
rect 24719 5556 24731 5559
rect 25038 5556 25044 5568
rect 24719 5528 25044 5556
rect 24719 5525 24731 5528
rect 24673 5519 24731 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 25133 5559 25191 5565
rect 25133 5525 25145 5559
rect 25179 5556 25191 5559
rect 31570 5556 31576 5568
rect 25179 5528 31576 5556
rect 25179 5525 25191 5528
rect 25133 5519 25191 5525
rect 31570 5516 31576 5528
rect 31628 5516 31634 5568
rect 31726 5556 31754 5596
rect 36998 5584 37004 5636
rect 37056 5584 37062 5636
rect 46293 5627 46351 5633
rect 46293 5593 46305 5627
rect 46339 5624 46351 5627
rect 49510 5624 49516 5636
rect 46339 5596 49516 5624
rect 46339 5593 46351 5596
rect 46293 5587 46351 5593
rect 49510 5584 49516 5596
rect 49568 5584 49574 5636
rect 49605 5627 49663 5633
rect 49605 5593 49617 5627
rect 49651 5624 49663 5627
rect 52362 5624 52368 5636
rect 49651 5596 52368 5624
rect 49651 5593 49663 5596
rect 49605 5587 49663 5593
rect 52362 5584 52368 5596
rect 52420 5584 52426 5636
rect 33318 5556 33324 5568
rect 31726 5528 33324 5556
rect 33318 5516 33324 5528
rect 33376 5516 33382 5568
rect 35713 5559 35771 5565
rect 35713 5525 35725 5559
rect 35759 5556 35771 5559
rect 35894 5556 35900 5568
rect 35759 5528 35900 5556
rect 35759 5525 35771 5528
rect 35713 5519 35771 5525
rect 35894 5516 35900 5528
rect 35952 5516 35958 5568
rect 41690 5516 41696 5568
rect 41748 5516 41754 5568
rect 45922 5516 45928 5568
rect 45980 5556 45986 5568
rect 47394 5556 47400 5568
rect 45980 5528 47400 5556
rect 45980 5516 45986 5528
rect 47394 5516 47400 5528
rect 47452 5516 47458 5568
rect 52546 5516 52552 5568
rect 52604 5556 52610 5568
rect 52748 5556 52776 5655
rect 52914 5652 52920 5704
rect 52972 5692 52978 5704
rect 53377 5695 53435 5701
rect 53377 5692 53389 5695
rect 52972 5664 53389 5692
rect 52972 5652 52978 5664
rect 53377 5661 53389 5664
rect 53423 5661 53435 5695
rect 53377 5655 53435 5661
rect 53834 5652 53840 5704
rect 53892 5692 53898 5704
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53892 5664 54125 5692
rect 53892 5652 53898 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 56321 5695 56379 5701
rect 56321 5661 56333 5695
rect 56367 5692 56379 5695
rect 56410 5692 56416 5704
rect 56367 5664 56416 5692
rect 56367 5661 56379 5664
rect 56321 5655 56379 5661
rect 56410 5652 56416 5664
rect 56468 5692 56474 5704
rect 59556 5701 59584 5732
rect 57977 5695 58035 5701
rect 57977 5692 57989 5695
rect 56468 5664 57989 5692
rect 56468 5652 56474 5664
rect 57977 5661 57989 5664
rect 58023 5692 58035 5695
rect 59541 5695 59599 5701
rect 59541 5692 59553 5695
rect 58023 5664 59553 5692
rect 58023 5661 58035 5664
rect 57977 5655 58035 5661
rect 59541 5661 59553 5664
rect 59587 5661 59599 5695
rect 59541 5655 59599 5661
rect 59725 5695 59783 5701
rect 59725 5661 59737 5695
rect 59771 5692 59783 5695
rect 60734 5692 60740 5704
rect 59771 5664 60740 5692
rect 59771 5661 59783 5664
rect 59725 5655 59783 5661
rect 60734 5652 60740 5664
rect 60792 5652 60798 5704
rect 61120 5636 61148 5732
rect 61654 5720 61660 5772
rect 61712 5720 61718 5772
rect 62574 5720 62580 5772
rect 62632 5760 62638 5772
rect 64156 5760 64184 5800
rect 67634 5788 67640 5800
rect 67692 5788 67698 5840
rect 62632 5732 64184 5760
rect 65061 5763 65119 5769
rect 62632 5720 62638 5732
rect 65061 5729 65073 5763
rect 65107 5760 65119 5763
rect 65978 5760 65984 5772
rect 65107 5732 65984 5760
rect 65107 5729 65119 5732
rect 65061 5723 65119 5729
rect 65978 5720 65984 5732
rect 66036 5720 66042 5772
rect 66162 5720 66168 5772
rect 66220 5720 66226 5772
rect 68462 5720 68468 5772
rect 68520 5720 68526 5772
rect 61473 5695 61531 5701
rect 61473 5686 61485 5695
rect 61304 5661 61485 5686
rect 61519 5661 61531 5695
rect 61304 5658 61531 5661
rect 53006 5584 53012 5636
rect 53064 5624 53070 5636
rect 60918 5624 60924 5636
rect 53064 5596 60924 5624
rect 53064 5584 53070 5596
rect 60918 5584 60924 5596
rect 60976 5584 60982 5636
rect 61102 5584 61108 5636
rect 61160 5624 61166 5636
rect 61304 5624 61332 5658
rect 61473 5655 61531 5658
rect 61160 5596 61332 5624
rect 61160 5584 61166 5596
rect 52604 5528 52776 5556
rect 53285 5559 53343 5565
rect 52604 5516 52610 5528
rect 53285 5525 53297 5559
rect 53331 5556 53343 5559
rect 54662 5556 54668 5568
rect 53331 5528 54668 5556
rect 53331 5525 53343 5528
rect 53285 5519 53343 5525
rect 54662 5516 54668 5528
rect 54720 5516 54726 5568
rect 54757 5559 54815 5565
rect 54757 5525 54769 5559
rect 54803 5556 54815 5559
rect 54846 5556 54852 5568
rect 54803 5528 54852 5556
rect 54803 5525 54815 5528
rect 54757 5519 54815 5525
rect 54846 5516 54852 5528
rect 54904 5516 54910 5568
rect 55582 5516 55588 5568
rect 55640 5556 55646 5568
rect 55861 5559 55919 5565
rect 55861 5556 55873 5559
rect 55640 5528 55873 5556
rect 55640 5516 55646 5528
rect 55861 5525 55873 5528
rect 55907 5525 55919 5559
rect 55861 5519 55919 5525
rect 56137 5559 56195 5565
rect 56137 5525 56149 5559
rect 56183 5556 56195 5559
rect 56226 5556 56232 5568
rect 56183 5528 56232 5556
rect 56183 5525 56195 5528
rect 56137 5519 56195 5525
rect 56226 5516 56232 5528
rect 56284 5516 56290 5568
rect 56318 5516 56324 5568
rect 56376 5556 56382 5568
rect 59630 5556 59636 5568
rect 56376 5528 59636 5556
rect 56376 5516 56382 5528
rect 59630 5516 59636 5528
rect 59688 5516 59694 5568
rect 61194 5516 61200 5568
rect 61252 5556 61258 5568
rect 61289 5559 61347 5565
rect 61289 5556 61301 5559
rect 61252 5528 61301 5556
rect 61252 5516 61258 5528
rect 61289 5525 61301 5528
rect 61335 5525 61347 5559
rect 61485 5556 61513 5655
rect 62942 5652 62948 5704
rect 63000 5652 63006 5704
rect 63129 5695 63187 5701
rect 63129 5661 63141 5695
rect 63175 5692 63187 5695
rect 64877 5695 64935 5701
rect 64877 5692 64889 5695
rect 63175 5664 64889 5692
rect 63175 5661 63187 5664
rect 63129 5655 63187 5661
rect 63236 5556 63264 5664
rect 64877 5661 64889 5664
rect 64923 5692 64935 5695
rect 66349 5695 66407 5701
rect 66349 5692 66361 5695
rect 64923 5664 66361 5692
rect 64923 5661 64935 5664
rect 64877 5655 64935 5661
rect 66349 5661 66361 5664
rect 66395 5692 66407 5695
rect 68281 5695 68339 5701
rect 68281 5692 68293 5695
rect 66395 5664 68293 5692
rect 66395 5661 66407 5664
rect 66349 5655 66407 5661
rect 68281 5661 68293 5664
rect 68327 5661 68339 5695
rect 68281 5655 68339 5661
rect 63586 5584 63592 5636
rect 63644 5624 63650 5636
rect 65334 5624 65340 5636
rect 63644 5596 65340 5624
rect 63644 5584 63650 5596
rect 65334 5584 65340 5596
rect 65392 5584 65398 5636
rect 61485 5528 63264 5556
rect 61289 5519 61347 5525
rect 63310 5516 63316 5568
rect 63368 5516 63374 5568
rect 64693 5559 64751 5565
rect 64693 5525 64705 5559
rect 64739 5556 64751 5559
rect 64782 5556 64788 5568
rect 64739 5528 64788 5556
rect 64739 5525 64751 5528
rect 64693 5519 64751 5525
rect 64782 5516 64788 5528
rect 64840 5516 64846 5568
rect 66438 5516 66444 5568
rect 66496 5556 66502 5568
rect 66533 5559 66591 5565
rect 66533 5556 66545 5559
rect 66496 5528 66545 5556
rect 66496 5516 66502 5528
rect 66533 5525 66545 5528
rect 66579 5525 66591 5559
rect 66533 5519 66591 5525
rect 68094 5516 68100 5568
rect 68152 5516 68158 5568
rect 1012 5466 74980 5488
rect 1012 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74980 5466
rect 1012 5392 74980 5414
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 63586 5352 63592 5364
rect 26660 5324 63592 5352
rect 26660 5312 26666 5324
rect 63586 5312 63592 5324
rect 63644 5312 63650 5364
rect 24412 5256 26556 5284
rect 23934 5176 23940 5228
rect 23992 5216 23998 5228
rect 24412 5225 24440 5256
rect 24397 5219 24455 5225
rect 24397 5216 24409 5219
rect 23992 5188 24409 5216
rect 23992 5176 23998 5188
rect 24397 5185 24409 5188
rect 24443 5185 24455 5219
rect 24397 5179 24455 5185
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 25590 5176 25596 5228
rect 25648 5216 25654 5228
rect 25958 5216 25964 5228
rect 25648 5188 25964 5216
rect 25648 5176 25654 5188
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 26068 5225 26096 5256
rect 26528 5225 26556 5256
rect 26786 5244 26792 5296
rect 26844 5284 26850 5296
rect 31202 5284 31208 5296
rect 26844 5256 31208 5284
rect 26844 5244 26850 5256
rect 31202 5244 31208 5256
rect 31260 5244 31266 5296
rect 46198 5284 46204 5296
rect 31312 5256 46204 5284
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 26421 5219 26479 5225
rect 26421 5185 26433 5219
rect 26467 5185 26479 5219
rect 26421 5179 26479 5185
rect 26513 5219 26571 5225
rect 26513 5185 26525 5219
rect 26559 5216 26571 5219
rect 27249 5219 27307 5225
rect 27249 5216 27261 5219
rect 26559 5188 27261 5216
rect 26559 5185 26571 5188
rect 26513 5179 26571 5185
rect 27249 5185 27261 5188
rect 27295 5216 27307 5219
rect 27295 5188 27660 5216
rect 27295 5185 27307 5188
rect 27249 5179 27307 5185
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5148 24271 5151
rect 24578 5148 24584 5160
rect 24259 5120 24584 5148
rect 24259 5117 24271 5120
rect 24213 5111 24271 5117
rect 24578 5108 24584 5120
rect 24636 5108 24642 5160
rect 25406 5108 25412 5160
rect 25464 5108 25470 5160
rect 25866 5108 25872 5160
rect 25924 5108 25930 5160
rect 26436 5148 26464 5179
rect 26602 5148 26608 5160
rect 26436 5120 26608 5148
rect 26602 5108 26608 5120
rect 26660 5108 26666 5160
rect 27065 5151 27123 5157
rect 27065 5117 27077 5151
rect 27111 5117 27123 5151
rect 27065 5111 27123 5117
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 24673 5083 24731 5089
rect 24673 5080 24685 5083
rect 23532 5052 24685 5080
rect 23532 5040 23538 5052
rect 24673 5049 24685 5052
rect 24719 5049 24731 5083
rect 24673 5043 24731 5049
rect 25777 5083 25835 5089
rect 25777 5049 25789 5083
rect 25823 5080 25835 5083
rect 26786 5080 26792 5092
rect 25823 5052 26792 5080
rect 25823 5049 25835 5052
rect 25777 5043 25835 5049
rect 26786 5040 26792 5052
rect 26844 5040 26850 5092
rect 27080 5080 27108 5111
rect 27522 5108 27528 5160
rect 27580 5108 27586 5160
rect 27632 5148 27660 5188
rect 27706 5176 27712 5228
rect 27764 5216 27770 5228
rect 28166 5216 28172 5228
rect 27764 5188 28172 5216
rect 27764 5176 27770 5188
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 28261 5219 28319 5225
rect 28261 5185 28273 5219
rect 28307 5185 28319 5219
rect 28261 5179 28319 5185
rect 27982 5148 27988 5160
rect 27632 5120 27988 5148
rect 27982 5108 27988 5120
rect 28040 5148 28046 5160
rect 28276 5148 28304 5179
rect 28442 5176 28448 5228
rect 28500 5176 28506 5228
rect 28885 5217 28943 5223
rect 28885 5214 28897 5217
rect 28828 5186 28897 5214
rect 28828 5148 28856 5186
rect 28885 5183 28897 5186
rect 28931 5214 28943 5217
rect 29104 5216 29408 5222
rect 29549 5219 29607 5225
rect 29549 5216 29561 5219
rect 29012 5214 29561 5216
rect 28931 5194 29561 5214
rect 28931 5188 29132 5194
rect 29380 5188 29561 5194
rect 28931 5186 29040 5188
rect 28931 5183 28943 5186
rect 28885 5177 28943 5183
rect 29549 5185 29561 5188
rect 29595 5185 29607 5219
rect 29549 5179 29607 5185
rect 28040 5120 28856 5148
rect 29089 5151 29147 5157
rect 28040 5108 28046 5120
rect 29089 5117 29101 5151
rect 29135 5117 29147 5151
rect 29564 5148 29592 5179
rect 29638 5176 29644 5228
rect 29696 5176 29702 5228
rect 30101 5219 30159 5225
rect 30101 5185 30113 5219
rect 30147 5216 30159 5219
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 30147 5188 30665 5216
rect 30147 5185 30159 5188
rect 30101 5179 30159 5185
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 30116 5148 30144 5179
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 29564 5120 30144 5148
rect 29089 5111 29147 5117
rect 28994 5080 29000 5092
rect 27080 5052 29000 5080
rect 28994 5040 29000 5052
rect 29052 5040 29058 5092
rect 29104 5080 29132 5111
rect 30282 5108 30288 5160
rect 30340 5108 30346 5160
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 31312 5148 31340 5256
rect 46198 5244 46204 5256
rect 46256 5244 46262 5296
rect 46474 5244 46480 5296
rect 46532 5284 46538 5296
rect 59078 5284 59084 5296
rect 46532 5256 59084 5284
rect 46532 5244 46538 5256
rect 59078 5244 59084 5256
rect 59136 5244 59142 5296
rect 61010 5244 61016 5296
rect 61068 5284 61074 5296
rect 62850 5284 62856 5296
rect 61068 5256 62856 5284
rect 61068 5244 61074 5256
rect 62850 5244 62856 5256
rect 62908 5244 62914 5296
rect 69658 5244 69664 5296
rect 69716 5284 69722 5296
rect 69716 5256 73568 5284
rect 69716 5244 69722 5256
rect 31386 5176 31392 5228
rect 31444 5216 31450 5228
rect 31444 5188 42932 5216
rect 31444 5176 31450 5188
rect 30432 5120 31340 5148
rect 30432 5108 30438 5120
rect 40402 5108 40408 5160
rect 40460 5108 40466 5160
rect 41046 5108 41052 5160
rect 41104 5108 41110 5160
rect 41506 5108 41512 5160
rect 41564 5108 41570 5160
rect 42904 5148 42932 5188
rect 42978 5176 42984 5228
rect 43036 5176 43042 5228
rect 44177 5219 44235 5225
rect 44177 5185 44189 5219
rect 44223 5216 44235 5219
rect 45922 5216 45928 5228
rect 44223 5188 45928 5216
rect 44223 5185 44235 5188
rect 44177 5179 44235 5185
rect 45922 5176 45928 5188
rect 45980 5176 45986 5228
rect 46290 5176 46296 5228
rect 46348 5176 46354 5228
rect 47213 5219 47271 5225
rect 47213 5185 47225 5219
rect 47259 5216 47271 5219
rect 47259 5188 51074 5216
rect 47259 5185 47271 5188
rect 47213 5179 47271 5185
rect 44082 5148 44088 5160
rect 42904 5120 44088 5148
rect 44082 5108 44088 5120
rect 44140 5108 44146 5160
rect 44545 5151 44603 5157
rect 44545 5117 44557 5151
rect 44591 5148 44603 5151
rect 44634 5148 44640 5160
rect 44591 5120 44640 5148
rect 44591 5117 44603 5120
rect 44545 5111 44603 5117
rect 44634 5108 44640 5120
rect 44692 5108 44698 5160
rect 45370 5108 45376 5160
rect 45428 5108 45434 5160
rect 46014 5108 46020 5160
rect 46072 5148 46078 5160
rect 46109 5151 46167 5157
rect 46109 5148 46121 5151
rect 46072 5120 46121 5148
rect 46072 5108 46078 5120
rect 46109 5117 46121 5120
rect 46155 5117 46167 5151
rect 46109 5111 46167 5117
rect 46382 5108 46388 5160
rect 46440 5148 46446 5160
rect 46569 5151 46627 5157
rect 46569 5148 46581 5151
rect 46440 5120 46581 5148
rect 46440 5108 46446 5120
rect 46569 5117 46581 5120
rect 46615 5117 46627 5151
rect 46569 5111 46627 5117
rect 47486 5108 47492 5160
rect 47544 5108 47550 5160
rect 48038 5108 48044 5160
rect 48096 5148 48102 5160
rect 48133 5151 48191 5157
rect 48133 5148 48145 5151
rect 48096 5120 48145 5148
rect 48096 5108 48102 5120
rect 48133 5117 48145 5120
rect 48179 5117 48191 5151
rect 48133 5111 48191 5117
rect 49142 5108 49148 5160
rect 49200 5108 49206 5160
rect 49786 5108 49792 5160
rect 49844 5108 49850 5160
rect 51046 5148 51074 5188
rect 52362 5176 52368 5228
rect 52420 5216 52426 5228
rect 53006 5216 53012 5228
rect 52420 5188 53012 5216
rect 52420 5176 52426 5188
rect 53006 5176 53012 5188
rect 53064 5176 53070 5228
rect 53098 5176 53104 5228
rect 53156 5176 53162 5228
rect 54570 5216 54576 5228
rect 53208 5188 54576 5216
rect 53208 5148 53236 5188
rect 54570 5176 54576 5188
rect 54628 5176 54634 5228
rect 54757 5219 54815 5225
rect 54757 5185 54769 5219
rect 54803 5185 54815 5219
rect 54757 5179 54815 5185
rect 51046 5120 53236 5148
rect 53282 5108 53288 5160
rect 53340 5108 53346 5160
rect 53374 5108 53380 5160
rect 53432 5148 53438 5160
rect 54772 5148 54800 5179
rect 54938 5176 54944 5228
rect 54996 5176 55002 5228
rect 55030 5176 55036 5228
rect 55088 5216 55094 5228
rect 55088 5188 57974 5216
rect 55088 5176 55094 5188
rect 56410 5148 56416 5160
rect 53432 5120 56416 5148
rect 53432 5108 53438 5120
rect 56410 5108 56416 5120
rect 56468 5108 56474 5160
rect 57946 5148 57974 5188
rect 61286 5176 61292 5228
rect 61344 5216 61350 5228
rect 73540 5225 73568 5256
rect 70213 5219 70271 5225
rect 70213 5216 70225 5219
rect 61344 5188 70225 5216
rect 61344 5176 61350 5188
rect 70213 5185 70225 5188
rect 70259 5216 70271 5219
rect 71685 5219 71743 5225
rect 71685 5216 71697 5219
rect 70259 5188 71697 5216
rect 70259 5185 70271 5188
rect 70213 5179 70271 5185
rect 71685 5185 71697 5188
rect 71731 5216 71743 5219
rect 73433 5219 73491 5225
rect 73433 5216 73445 5219
rect 71731 5188 73445 5216
rect 71731 5185 71743 5188
rect 71685 5179 71743 5185
rect 73433 5185 73445 5188
rect 73479 5185 73491 5219
rect 73433 5179 73491 5185
rect 73525 5219 73583 5225
rect 73525 5185 73537 5219
rect 73571 5185 73583 5219
rect 73525 5179 73583 5185
rect 65426 5148 65432 5160
rect 57946 5120 65432 5148
rect 65426 5108 65432 5120
rect 65484 5108 65490 5160
rect 69934 5108 69940 5160
rect 69992 5148 69998 5160
rect 70397 5151 70455 5157
rect 70397 5148 70409 5151
rect 69992 5120 70409 5148
rect 69992 5108 69998 5120
rect 70397 5117 70409 5120
rect 70443 5117 70455 5151
rect 70397 5111 70455 5117
rect 71869 5151 71927 5157
rect 71869 5117 71881 5151
rect 71915 5117 71927 5151
rect 71869 5111 71927 5117
rect 29270 5080 29276 5092
rect 29104 5052 29276 5080
rect 29270 5040 29276 5052
rect 29328 5040 29334 5092
rect 29638 5040 29644 5092
rect 29696 5080 29702 5092
rect 47026 5080 47032 5092
rect 29696 5052 46244 5080
rect 29696 5040 29702 5052
rect 24581 5015 24639 5021
rect 24581 4981 24593 5015
rect 24627 5012 24639 5015
rect 26142 5012 26148 5024
rect 24627 4984 26148 5012
rect 24627 4981 24639 4984
rect 24581 4975 24639 4981
rect 26142 4972 26148 4984
rect 26200 4972 26206 5024
rect 26234 4972 26240 5024
rect 26292 4972 26298 5024
rect 26694 4972 26700 5024
rect 26752 4972 26758 5024
rect 27433 5015 27491 5021
rect 27433 4981 27445 5015
rect 27479 5012 27491 5015
rect 27798 5012 27804 5024
rect 27479 4984 27804 5012
rect 27479 4981 27491 4984
rect 27433 4975 27491 4981
rect 27798 4972 27804 4984
rect 27856 4972 27862 5024
rect 27890 4972 27896 5024
rect 27948 4972 27954 5024
rect 28077 5015 28135 5021
rect 28077 4981 28089 5015
rect 28123 5012 28135 5015
rect 28534 5012 28540 5024
rect 28123 4984 28540 5012
rect 28123 4981 28135 4984
rect 28077 4975 28135 4981
rect 28534 4972 28540 4984
rect 28592 4972 28598 5024
rect 28718 4972 28724 5024
rect 28776 4972 28782 5024
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 29086 5012 29092 5024
rect 28868 4984 29092 5012
rect 28868 4972 28874 4984
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 29362 4972 29368 5024
rect 29420 4972 29426 5024
rect 29454 4972 29460 5024
rect 29512 5012 29518 5024
rect 29917 5015 29975 5021
rect 29917 5012 29929 5015
rect 29512 4984 29929 5012
rect 29512 4972 29518 4984
rect 29917 4981 29929 4984
rect 29963 4981 29975 5015
rect 29917 4975 29975 4981
rect 30466 4972 30472 5024
rect 30524 4972 30530 5024
rect 42153 5015 42211 5021
rect 42153 4981 42165 5015
rect 42199 5012 42211 5015
rect 45002 5012 45008 5024
rect 42199 4984 45008 5012
rect 42199 4981 42211 4984
rect 42153 4975 42211 4981
rect 45002 4972 45008 4984
rect 45060 4972 45066 5024
rect 45094 4972 45100 5024
rect 45152 4972 45158 5024
rect 46017 5015 46075 5021
rect 46017 4981 46029 5015
rect 46063 5012 46075 5015
rect 46106 5012 46112 5024
rect 46063 4984 46112 5012
rect 46063 4981 46075 4984
rect 46017 4975 46075 4981
rect 46106 4972 46112 4984
rect 46164 4972 46170 5024
rect 46216 5012 46244 5052
rect 46400 5052 47032 5080
rect 46400 5012 46428 5052
rect 47026 5040 47032 5052
rect 47084 5040 47090 5092
rect 47302 5040 47308 5092
rect 47360 5080 47366 5092
rect 63770 5080 63776 5092
rect 47360 5052 63776 5080
rect 47360 5040 47366 5052
rect 63770 5040 63776 5052
rect 63828 5040 63834 5092
rect 69750 5040 69756 5092
rect 69808 5080 69814 5092
rect 71884 5080 71912 5111
rect 69808 5052 71912 5080
rect 69808 5040 69814 5052
rect 46216 4984 46428 5012
rect 46477 5015 46535 5021
rect 46477 4981 46489 5015
rect 46523 5012 46535 5015
rect 47118 5012 47124 5024
rect 46523 4984 47124 5012
rect 46523 4981 46535 4984
rect 46477 4975 46535 4981
rect 47118 4972 47124 4984
rect 47176 4972 47182 5024
rect 47394 4972 47400 5024
rect 47452 5012 47458 5024
rect 49326 5012 49332 5024
rect 47452 4984 49332 5012
rect 47452 4972 47458 4984
rect 49326 4972 49332 4984
rect 49384 4972 49390 5024
rect 52914 4972 52920 5024
rect 52972 4972 52978 5024
rect 54573 5015 54631 5021
rect 54573 4981 54585 5015
rect 54619 5012 54631 5015
rect 54662 5012 54668 5024
rect 54619 4984 54668 5012
rect 54619 4981 54631 4984
rect 54573 4975 54631 4981
rect 54662 4972 54668 4984
rect 54720 4972 54726 5024
rect 54754 4972 54760 5024
rect 54812 5012 54818 5024
rect 63494 5012 63500 5024
rect 54812 4984 63500 5012
rect 54812 4972 54818 4984
rect 63494 4972 63500 4984
rect 63552 4972 63558 5024
rect 69842 4972 69848 5024
rect 69900 5012 69906 5024
rect 70029 5015 70087 5021
rect 70029 5012 70041 5015
rect 69900 4984 70041 5012
rect 69900 4972 69906 4984
rect 70029 4981 70041 4984
rect 70075 4981 70087 5015
rect 70029 4975 70087 4981
rect 71406 4972 71412 5024
rect 71464 5012 71470 5024
rect 71501 5015 71559 5021
rect 71501 5012 71513 5015
rect 71464 4984 71513 5012
rect 71464 4972 71470 4984
rect 71501 4981 71513 4984
rect 71547 4981 71559 5015
rect 71501 4975 71559 4981
rect 73246 4972 73252 5024
rect 73304 4972 73310 5024
rect 1012 4922 74980 4944
rect 1012 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 74980 4922
rect 1012 4848 74980 4870
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 30006 4808 30012 4820
rect 26292 4780 30012 4808
rect 26292 4768 26298 4780
rect 30006 4768 30012 4780
rect 30064 4768 30070 4820
rect 32306 4768 32312 4820
rect 32364 4808 32370 4820
rect 41506 4808 41512 4820
rect 32364 4780 41512 4808
rect 32364 4768 32370 4780
rect 41506 4768 41512 4780
rect 41564 4768 41570 4820
rect 42610 4768 42616 4820
rect 42668 4768 42674 4820
rect 45094 4768 45100 4820
rect 45152 4808 45158 4820
rect 61010 4808 61016 4820
rect 45152 4780 61016 4808
rect 45152 4768 45158 4780
rect 61010 4768 61016 4780
rect 61068 4768 61074 4820
rect 62758 4768 62764 4820
rect 62816 4808 62822 4820
rect 68738 4808 68744 4820
rect 62816 4780 68744 4808
rect 62816 4768 62822 4780
rect 68738 4768 68744 4780
rect 68796 4768 68802 4820
rect 25590 4700 25596 4752
rect 25648 4740 25654 4752
rect 27706 4740 27712 4752
rect 25648 4712 27712 4740
rect 25648 4700 25654 4712
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 27890 4700 27896 4752
rect 27948 4740 27954 4752
rect 27948 4712 34284 4740
rect 27948 4700 27954 4712
rect 24578 4632 24584 4684
rect 24636 4672 24642 4684
rect 31386 4672 31392 4684
rect 24636 4644 31392 4672
rect 24636 4632 24642 4644
rect 31386 4632 31392 4644
rect 31444 4632 31450 4684
rect 34054 4632 34060 4684
rect 34112 4672 34118 4684
rect 34149 4675 34207 4681
rect 34149 4672 34161 4675
rect 34112 4644 34161 4672
rect 34112 4632 34118 4644
rect 34149 4641 34161 4644
rect 34195 4641 34207 4675
rect 34256 4672 34284 4712
rect 35066 4700 35072 4752
rect 35124 4740 35130 4752
rect 42978 4740 42984 4752
rect 35124 4712 42984 4740
rect 35124 4700 35130 4712
rect 42978 4700 42984 4712
rect 43036 4700 43042 4752
rect 44726 4740 44732 4752
rect 44100 4712 44732 4740
rect 36814 4672 36820 4684
rect 34256 4644 36820 4672
rect 34149 4635 34207 4641
rect 36814 4632 36820 4644
rect 36872 4632 36878 4684
rect 44100 4681 44128 4712
rect 44726 4700 44732 4712
rect 44784 4700 44790 4752
rect 45002 4700 45008 4752
rect 45060 4740 45066 4752
rect 45060 4712 49280 4740
rect 45060 4700 45066 4712
rect 44085 4675 44143 4681
rect 44085 4641 44097 4675
rect 44131 4641 44143 4675
rect 44085 4635 44143 4641
rect 46308 4644 46888 4672
rect 46308 4616 46336 4644
rect 26694 4564 26700 4616
rect 26752 4604 26758 4616
rect 28994 4604 29000 4616
rect 26752 4576 29000 4604
rect 26752 4564 26758 4576
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 29086 4564 29092 4616
rect 29144 4604 29150 4616
rect 29144 4576 31754 4604
rect 29144 4564 29150 4576
rect 25406 4496 25412 4548
rect 25464 4536 25470 4548
rect 30098 4536 30104 4548
rect 25464 4508 30104 4536
rect 25464 4496 25470 4508
rect 30098 4496 30104 4508
rect 30156 4496 30162 4548
rect 26142 4428 26148 4480
rect 26200 4468 26206 4480
rect 29638 4468 29644 4480
rect 26200 4440 29644 4468
rect 26200 4428 26206 4440
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 31726 4468 31754 4576
rect 33962 4564 33968 4616
rect 34020 4564 34026 4616
rect 41230 4564 41236 4616
rect 41288 4564 41294 4616
rect 41690 4564 41696 4616
rect 41748 4604 41754 4616
rect 41969 4607 42027 4613
rect 41969 4604 41981 4607
rect 41748 4576 41981 4604
rect 41748 4564 41754 4576
rect 41969 4573 41981 4576
rect 42015 4573 42027 4607
rect 41969 4567 42027 4573
rect 43346 4564 43352 4616
rect 43404 4564 43410 4616
rect 44269 4607 44327 4613
rect 44269 4604 44281 4607
rect 44192 4598 44281 4604
rect 44100 4576 44281 4598
rect 44100 4570 44220 4576
rect 44269 4573 44281 4576
rect 44315 4604 44327 4607
rect 46290 4604 46296 4616
rect 44315 4576 46296 4604
rect 44315 4573 44327 4576
rect 32582 4496 32588 4548
rect 32640 4536 32646 4548
rect 36538 4536 36544 4548
rect 32640 4508 36544 4536
rect 32640 4496 32646 4508
rect 36538 4496 36544 4508
rect 36596 4496 36602 4548
rect 44100 4536 44128 4570
rect 44269 4567 44327 4573
rect 46290 4564 46296 4576
rect 46348 4564 46354 4616
rect 46658 4564 46664 4616
rect 46716 4564 46722 4616
rect 46860 4615 46888 4644
rect 47026 4632 47032 4684
rect 47084 4672 47090 4684
rect 49252 4672 49280 4712
rect 49326 4700 49332 4752
rect 49384 4740 49390 4752
rect 65150 4740 65156 4752
rect 49384 4712 65156 4740
rect 49384 4700 49390 4712
rect 65150 4700 65156 4712
rect 65208 4700 65214 4752
rect 47084 4644 49188 4672
rect 49252 4644 51074 4672
rect 47084 4632 47090 4644
rect 46831 4609 46889 4615
rect 46831 4575 46843 4609
rect 46877 4575 46889 4609
rect 46831 4569 46889 4575
rect 46566 4536 46572 4548
rect 38626 4508 44128 4536
rect 44376 4508 46572 4536
rect 34698 4468 34704 4480
rect 31726 4440 34704 4468
rect 34698 4428 34704 4440
rect 34756 4468 34762 4480
rect 38626 4468 38654 4508
rect 34756 4440 38654 4468
rect 41877 4471 41935 4477
rect 34756 4428 34762 4440
rect 41877 4437 41889 4471
rect 41923 4468 41935 4471
rect 43898 4468 43904 4480
rect 41923 4440 43904 4468
rect 41923 4437 41935 4440
rect 41877 4431 41935 4437
rect 43898 4428 43904 4440
rect 43956 4428 43962 4480
rect 43993 4471 44051 4477
rect 43993 4437 44005 4471
rect 44039 4468 44051 4471
rect 44376 4468 44404 4508
rect 46566 4496 46572 4508
rect 46624 4496 46630 4548
rect 48958 4536 48964 4548
rect 46952 4508 48964 4536
rect 44039 4440 44404 4468
rect 44453 4471 44511 4477
rect 44039 4437 44051 4440
rect 43993 4431 44051 4437
rect 44453 4437 44465 4471
rect 44499 4468 44511 4471
rect 45922 4468 45928 4480
rect 44499 4440 45928 4468
rect 44499 4437 44511 4440
rect 44453 4431 44511 4437
rect 45922 4428 45928 4440
rect 45980 4428 45986 4480
rect 46750 4428 46756 4480
rect 46808 4468 46814 4480
rect 46952 4468 46980 4508
rect 48958 4496 48964 4508
rect 49016 4496 49022 4548
rect 49160 4536 49188 4644
rect 51046 4604 51074 4644
rect 51534 4632 51540 4684
rect 51592 4672 51598 4684
rect 54846 4672 54852 4684
rect 51592 4644 54852 4672
rect 51592 4632 51598 4644
rect 54846 4632 54852 4644
rect 54904 4632 54910 4684
rect 54938 4632 54944 4684
rect 54996 4672 55002 4684
rect 70762 4672 70768 4684
rect 54996 4644 70768 4672
rect 54996 4632 55002 4644
rect 70762 4632 70768 4644
rect 70820 4632 70826 4684
rect 61010 4604 61016 4616
rect 51046 4576 61016 4604
rect 61010 4564 61016 4576
rect 61068 4564 61074 4616
rect 61197 4607 61255 4613
rect 61197 4573 61209 4607
rect 61243 4604 61255 4607
rect 61286 4604 61292 4616
rect 61243 4576 61292 4604
rect 61243 4573 61255 4576
rect 61197 4567 61255 4573
rect 61286 4564 61292 4576
rect 61344 4564 61350 4616
rect 61470 4564 61476 4616
rect 61528 4604 61534 4616
rect 68554 4604 68560 4616
rect 61528 4576 68560 4604
rect 61528 4564 61534 4576
rect 68554 4564 68560 4576
rect 68612 4564 68618 4616
rect 60918 4536 60924 4548
rect 49160 4508 60924 4536
rect 60918 4496 60924 4508
rect 60976 4496 60982 4548
rect 61028 4508 61240 4536
rect 46808 4440 46980 4468
rect 47029 4471 47087 4477
rect 46808 4428 46814 4440
rect 47029 4437 47041 4471
rect 47075 4468 47087 4471
rect 49050 4468 49056 4480
rect 47075 4440 49056 4468
rect 47075 4437 47087 4440
rect 47029 4431 47087 4437
rect 49050 4428 49056 4440
rect 49108 4428 49114 4480
rect 55490 4428 55496 4480
rect 55548 4468 55554 4480
rect 61028 4468 61056 4508
rect 55548 4440 61056 4468
rect 55548 4428 55554 4440
rect 61102 4428 61108 4480
rect 61160 4428 61166 4480
rect 61212 4468 61240 4508
rect 62850 4496 62856 4548
rect 62908 4536 62914 4548
rect 69290 4536 69296 4548
rect 62908 4508 69296 4536
rect 62908 4496 62914 4508
rect 69290 4496 69296 4508
rect 69348 4496 69354 4548
rect 68002 4468 68008 4480
rect 61212 4440 68008 4468
rect 68002 4428 68008 4440
rect 68060 4428 68066 4480
rect 1012 4378 74980 4400
rect 1012 4326 4210 4378
rect 4262 4326 4274 4378
rect 4326 4326 4338 4378
rect 4390 4326 4402 4378
rect 4454 4326 4466 4378
rect 4518 4326 14210 4378
rect 14262 4326 14274 4378
rect 14326 4326 14338 4378
rect 14390 4326 14402 4378
rect 14454 4326 14466 4378
rect 14518 4326 24210 4378
rect 24262 4326 24274 4378
rect 24326 4326 24338 4378
rect 24390 4326 24402 4378
rect 24454 4326 24466 4378
rect 24518 4326 34210 4378
rect 34262 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 44210 4378
rect 44262 4326 44274 4378
rect 44326 4326 44338 4378
rect 44390 4326 44402 4378
rect 44454 4326 44466 4378
rect 44518 4326 54210 4378
rect 54262 4326 54274 4378
rect 54326 4326 54338 4378
rect 54390 4326 54402 4378
rect 54454 4326 54466 4378
rect 54518 4326 64210 4378
rect 64262 4326 64274 4378
rect 64326 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 74210 4378
rect 74262 4326 74274 4378
rect 74326 4326 74338 4378
rect 74390 4326 74402 4378
rect 74454 4326 74466 4378
rect 74518 4326 74980 4378
rect 1012 4304 74980 4326
rect 27614 4224 27620 4276
rect 27672 4264 27678 4276
rect 34790 4264 34796 4276
rect 27672 4236 34796 4264
rect 27672 4224 27678 4236
rect 34790 4224 34796 4236
rect 34848 4224 34854 4276
rect 36538 4224 36544 4276
rect 36596 4264 36602 4276
rect 47486 4264 47492 4276
rect 36596 4236 47492 4264
rect 36596 4224 36602 4236
rect 47486 4224 47492 4236
rect 47544 4224 47550 4276
rect 47578 4224 47584 4276
rect 47636 4264 47642 4276
rect 51534 4264 51540 4276
rect 47636 4236 51540 4264
rect 47636 4224 47642 4236
rect 51534 4224 51540 4236
rect 51592 4224 51598 4276
rect 53282 4224 53288 4276
rect 53340 4264 53346 4276
rect 62666 4264 62672 4276
rect 53340 4236 62672 4264
rect 53340 4224 53346 4236
rect 62666 4224 62672 4236
rect 62724 4224 62730 4276
rect 19628 4168 20392 4196
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 19628 4128 19656 4168
rect 19116 4100 19656 4128
rect 19705 4131 19763 4137
rect 19116 4088 19122 4100
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 20254 4128 20260 4140
rect 19751 4100 20260 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20364 4128 20392 4168
rect 27540 4168 29960 4196
rect 27540 4128 27568 4168
rect 20364 4100 27568 4128
rect 27614 4088 27620 4140
rect 27672 4088 27678 4140
rect 29932 4128 29960 4168
rect 30098 4156 30104 4208
rect 30156 4196 30162 4208
rect 65518 4196 65524 4208
rect 30156 4168 47440 4196
rect 30156 4156 30162 4168
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 27724 4100 29868 4128
rect 29932 4100 30849 4128
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 27724 4060 27752 4100
rect 19567 4032 27752 4060
rect 27893 4063 27951 4069
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 27893 4029 27905 4063
rect 27939 4060 27951 4063
rect 27982 4060 27988 4072
rect 27939 4032 27988 4060
rect 27939 4029 27951 4032
rect 27893 4023 27951 4029
rect 27982 4020 27988 4032
rect 28040 4020 28046 4072
rect 29730 4020 29736 4072
rect 29788 4020 29794 4072
rect 29840 4060 29868 4100
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 34606 4128 34612 4140
rect 31536 4100 34612 4128
rect 31536 4088 31542 4100
rect 34606 4088 34612 4100
rect 34664 4088 34670 4140
rect 34698 4088 34704 4140
rect 34756 4088 34762 4140
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 34885 4131 34943 4137
rect 34885 4128 34897 4131
rect 34848 4100 34897 4128
rect 34848 4088 34854 4100
rect 34885 4097 34897 4100
rect 34931 4097 34943 4131
rect 34885 4091 34943 4097
rect 34974 4088 34980 4140
rect 35032 4128 35038 4140
rect 42978 4128 42984 4140
rect 35032 4100 42984 4128
rect 35032 4088 35038 4100
rect 42978 4088 42984 4100
rect 43036 4088 43042 4140
rect 43898 4088 43904 4140
rect 43956 4128 43962 4140
rect 47026 4128 47032 4140
rect 43956 4100 47032 4128
rect 43956 4088 43962 4100
rect 47026 4088 47032 4100
rect 47084 4088 47090 4140
rect 47412 4128 47440 4168
rect 47688 4168 65524 4196
rect 47688 4128 47716 4168
rect 65518 4156 65524 4168
rect 65576 4156 65582 4208
rect 47412 4100 47716 4128
rect 48958 4088 48964 4140
rect 49016 4128 49022 4140
rect 55490 4128 55496 4140
rect 49016 4100 55496 4128
rect 49016 4088 49022 4100
rect 55490 4088 55496 4100
rect 55548 4088 55554 4140
rect 60734 4088 60740 4140
rect 60792 4128 60798 4140
rect 66622 4128 66628 4140
rect 60792 4100 66628 4128
rect 60792 4088 60798 4100
rect 66622 4088 66628 4100
rect 66680 4088 66686 4140
rect 41690 4060 41696 4072
rect 29840 4032 41696 4060
rect 41690 4020 41696 4032
rect 41748 4020 41754 4072
rect 61470 4020 61476 4072
rect 61528 4060 61534 4072
rect 66530 4060 66536 4072
rect 61528 4032 66536 4060
rect 61528 4020 61534 4032
rect 66530 4020 66536 4032
rect 66588 4020 66594 4072
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 40402 3992 40408 4004
rect 17920 3964 40408 3992
rect 17920 3952 17926 3964
rect 40402 3952 40408 3964
rect 40460 3952 40466 4004
rect 47026 3952 47032 4004
rect 47084 3992 47090 4004
rect 51258 3992 51264 4004
rect 47084 3964 51264 3992
rect 47084 3952 47090 3964
rect 51258 3952 51264 3964
rect 51316 3952 51322 4004
rect 60918 3952 60924 4004
rect 60976 3992 60982 4004
rect 62758 3992 62764 4004
rect 60976 3964 62764 3992
rect 60976 3952 60982 3964
rect 62758 3952 62764 3964
rect 62816 3952 62822 4004
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 27614 3924 27620 3936
rect 23440 3896 27620 3924
rect 23440 3884 23446 3896
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 30377 3927 30435 3933
rect 30377 3893 30389 3927
rect 30423 3924 30435 3927
rect 33962 3924 33968 3936
rect 30423 3896 33968 3924
rect 30423 3893 30435 3896
rect 30377 3887 30435 3893
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 35802 3924 35808 3936
rect 34848 3896 35808 3924
rect 34848 3884 34854 3896
rect 35802 3884 35808 3896
rect 35860 3884 35866 3936
rect 36998 3884 37004 3936
rect 37056 3924 37062 3936
rect 47394 3924 47400 3936
rect 37056 3896 47400 3924
rect 37056 3884 37062 3896
rect 47394 3884 47400 3896
rect 47452 3884 47458 3936
rect 1012 3834 74980 3856
rect 1012 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 74980 3834
rect 1012 3760 74980 3782
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 25590 3720 25596 3732
rect 20956 3692 25596 3720
rect 20956 3680 20962 3692
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 26050 3680 26056 3732
rect 26108 3680 26114 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 29730 3720 29736 3732
rect 26283 3692 29736 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 29730 3680 29736 3692
rect 29788 3680 29794 3732
rect 32306 3720 32312 3732
rect 31726 3692 32312 3720
rect 25774 3652 25780 3664
rect 19444 3624 25780 3652
rect 19444 3593 19472 3624
rect 25774 3612 25780 3624
rect 25832 3612 25838 3664
rect 31726 3652 31754 3692
rect 32306 3680 32312 3692
rect 32364 3680 32370 3732
rect 33045 3723 33103 3729
rect 33045 3689 33057 3723
rect 33091 3720 33103 3723
rect 33091 3692 33180 3720
rect 33091 3689 33103 3692
rect 33045 3683 33103 3689
rect 26896 3624 31754 3652
rect 31849 3655 31907 3661
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3553 19487 3587
rect 19429 3547 19487 3553
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3584 20039 3587
rect 26896 3584 26924 3624
rect 31849 3621 31861 3655
rect 31895 3652 31907 3655
rect 32674 3652 32680 3664
rect 31895 3624 32680 3652
rect 31895 3621 31907 3624
rect 31849 3615 31907 3621
rect 32674 3612 32680 3624
rect 32732 3612 32738 3664
rect 27890 3584 27896 3596
rect 20027 3556 26924 3584
rect 26988 3556 27896 3584
rect 20027 3553 20039 3556
rect 19981 3547 20039 3553
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19153 3519 19211 3525
rect 19153 3516 19165 3519
rect 18288 3488 19165 3516
rect 18288 3476 18294 3488
rect 19153 3485 19165 3488
rect 19199 3485 19211 3519
rect 19153 3479 19211 3485
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20530 3516 20536 3528
rect 20211 3488 20536 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22520 3488 22569 3516
rect 22520 3476 22526 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23440 3488 23489 3516
rect 23440 3476 23446 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 23584 3448 23612 3479
rect 24946 3476 24952 3528
rect 25004 3476 25010 3528
rect 25222 3476 25228 3528
rect 25280 3476 25286 3528
rect 25498 3476 25504 3528
rect 25556 3476 25562 3528
rect 25774 3476 25780 3528
rect 25832 3476 25838 3528
rect 25958 3476 25964 3528
rect 26016 3516 26022 3528
rect 26988 3516 27016 3556
rect 27890 3544 27896 3556
rect 27948 3544 27954 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 32766 3584 32772 3596
rect 28224 3556 32772 3584
rect 28224 3544 28230 3556
rect 32766 3544 32772 3556
rect 32824 3544 32830 3596
rect 33152 3584 33180 3692
rect 33226 3680 33232 3732
rect 33284 3720 33290 3732
rect 41230 3720 41236 3732
rect 33284 3692 41236 3720
rect 33284 3680 33290 3692
rect 41230 3680 41236 3692
rect 41288 3680 41294 3732
rect 36170 3612 36176 3664
rect 36228 3652 36234 3664
rect 49142 3652 49148 3664
rect 36228 3624 49148 3652
rect 36228 3612 36234 3624
rect 49142 3612 49148 3624
rect 49200 3612 49206 3664
rect 33152 3556 35940 3584
rect 26016 3488 27016 3516
rect 28077 3519 28135 3525
rect 26016 3476 26022 3488
rect 28077 3485 28089 3519
rect 28123 3516 28135 3519
rect 28718 3516 28724 3528
rect 28123 3488 28724 3516
rect 28123 3485 28135 3488
rect 28077 3479 28135 3485
rect 28718 3476 28724 3488
rect 28776 3476 28782 3528
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 31570 3476 31576 3528
rect 31628 3516 31634 3528
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31628 3488 31677 3516
rect 31628 3476 31634 3488
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 32214 3476 32220 3528
rect 32272 3476 32278 3528
rect 32858 3476 32864 3528
rect 32916 3476 32922 3528
rect 35912 3516 35940 3556
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 44634 3584 44640 3596
rect 36136 3556 44640 3584
rect 36136 3544 36142 3556
rect 44634 3544 44640 3556
rect 44692 3544 44698 3596
rect 52546 3584 52552 3596
rect 48286 3556 52552 3584
rect 37090 3516 37096 3528
rect 32968 3488 33180 3516
rect 35912 3488 37096 3516
rect 22066 3420 23612 3448
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 22066 3380 22094 3420
rect 25590 3408 25596 3460
rect 25648 3448 25654 3460
rect 25869 3451 25927 3457
rect 25869 3448 25881 3451
rect 25648 3420 25881 3448
rect 25648 3408 25654 3420
rect 25869 3417 25881 3420
rect 25915 3417 25927 3451
rect 25869 3411 25927 3417
rect 27706 3408 27712 3460
rect 27764 3408 27770 3460
rect 32968 3448 32996 3488
rect 27816 3420 32996 3448
rect 33152 3448 33180 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 42242 3476 42248 3528
rect 42300 3516 42306 3528
rect 48286 3516 48314 3556
rect 52546 3544 52552 3556
rect 52604 3544 52610 3596
rect 55858 3544 55864 3596
rect 55916 3584 55922 3596
rect 66346 3584 66352 3596
rect 55916 3556 66352 3584
rect 55916 3544 55922 3556
rect 66346 3544 66352 3556
rect 66404 3544 66410 3596
rect 42300 3488 48314 3516
rect 42300 3476 42306 3488
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 67358 3516 67364 3528
rect 51224 3488 67364 3516
rect 51224 3476 51230 3488
rect 67358 3476 67364 3488
rect 67416 3476 67422 3528
rect 45370 3448 45376 3460
rect 33152 3420 45376 3448
rect 20680 3352 22094 3380
rect 20680 3340 20686 3352
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 23201 3383 23259 3389
rect 23201 3380 23213 3383
rect 23164 3352 23213 3380
rect 23164 3340 23170 3352
rect 23201 3349 23213 3352
rect 23247 3349 23259 3383
rect 23201 3343 23259 3349
rect 23290 3340 23296 3392
rect 23348 3340 23354 3392
rect 26074 3383 26132 3389
rect 26074 3349 26086 3383
rect 26120 3380 26132 3383
rect 26234 3380 26240 3392
rect 26120 3352 26240 3380
rect 26120 3349 26132 3352
rect 26074 3343 26132 3349
rect 26234 3340 26240 3352
rect 26292 3380 26298 3392
rect 27154 3380 27160 3392
rect 26292 3352 27160 3380
rect 26292 3340 26298 3352
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 27617 3383 27675 3389
rect 27617 3349 27629 3383
rect 27663 3380 27675 3383
rect 27816 3380 27844 3420
rect 45370 3408 45376 3420
rect 45428 3408 45434 3460
rect 61378 3448 61384 3460
rect 51046 3420 61384 3448
rect 27663 3352 27844 3380
rect 27663 3349 27675 3352
rect 27617 3343 27675 3349
rect 27890 3340 27896 3392
rect 27948 3340 27954 3392
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 31294 3380 31300 3392
rect 28040 3352 31300 3380
rect 28040 3340 28046 3352
rect 31294 3340 31300 3352
rect 31352 3340 31358 3392
rect 31386 3340 31392 3392
rect 31444 3340 31450 3392
rect 32401 3383 32459 3389
rect 32401 3349 32413 3383
rect 32447 3380 32459 3383
rect 39758 3380 39764 3392
rect 32447 3352 39764 3380
rect 32447 3349 32459 3352
rect 32401 3343 32459 3349
rect 39758 3340 39764 3352
rect 39816 3340 39822 3392
rect 44910 3340 44916 3392
rect 44968 3380 44974 3392
rect 51046 3380 51074 3420
rect 61378 3408 61384 3420
rect 61436 3408 61442 3460
rect 44968 3352 51074 3380
rect 44968 3340 44974 3352
rect 1012 3290 74980 3312
rect 1012 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74980 3290
rect 1012 3216 74980 3238
rect 20530 3136 20536 3188
rect 20588 3136 20594 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 24854 3176 24860 3188
rect 21315 3148 24860 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 25774 3136 25780 3188
rect 25832 3176 25838 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25832 3148 25881 3176
rect 25832 3136 25838 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 27706 3136 27712 3188
rect 27764 3176 27770 3188
rect 28077 3179 28135 3185
rect 28077 3176 28089 3179
rect 27764 3148 28089 3176
rect 27764 3136 27770 3148
rect 28077 3145 28089 3148
rect 28123 3145 28135 3179
rect 28077 3139 28135 3145
rect 29457 3179 29515 3185
rect 29457 3145 29469 3179
rect 29503 3176 29515 3179
rect 29546 3176 29552 3188
rect 29503 3148 29552 3176
rect 29503 3145 29515 3148
rect 29457 3139 29515 3145
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 30193 3179 30251 3185
rect 30193 3145 30205 3179
rect 30239 3145 30251 3179
rect 33226 3176 33232 3188
rect 30193 3139 30251 3145
rect 32508 3148 33232 3176
rect 17862 3068 17868 3120
rect 17920 3068 17926 3120
rect 21110 3111 21168 3117
rect 21110 3077 21122 3111
rect 21156 3108 21168 3111
rect 21156 3080 22876 3108
rect 21156 3077 21168 3080
rect 21110 3071 21168 3077
rect 18138 3000 18144 3052
rect 18196 3000 18202 3052
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 20772 3012 21373 3040
rect 20772 3000 20778 3012
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 22738 3040 22744 3052
rect 21361 3003 21419 3009
rect 21468 3012 22744 3040
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 18969 2975 19027 2981
rect 18969 2972 18981 2975
rect 18748 2944 18981 2972
rect 18748 2932 18754 2944
rect 18969 2941 18981 2944
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 19150 2932 19156 2984
rect 19208 2932 19214 2984
rect 19886 2932 19892 2984
rect 19944 2932 19950 2984
rect 20898 2932 20904 2984
rect 20956 2932 20962 2984
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2972 21051 2975
rect 21468 2972 21496 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 21039 2944 21496 2972
rect 21039 2941 21051 2944
rect 20993 2935 21051 2941
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 21008 2904 21036 2935
rect 21726 2932 21732 2984
rect 21784 2932 21790 2984
rect 20588 2876 21036 2904
rect 20588 2864 20594 2876
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 22336 2876 22477 2904
rect 22336 2864 22342 2876
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22848 2904 22876 3080
rect 22922 3068 22928 3120
rect 22980 3108 22986 3120
rect 26050 3108 26056 3120
rect 22980 3080 26056 3108
rect 22980 3068 22986 3080
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 29362 3108 29368 3120
rect 26712 3080 29368 3108
rect 23106 3000 23112 3052
rect 23164 3000 23170 3052
rect 26712 3049 26740 3080
rect 29362 3068 29368 3080
rect 29420 3068 29426 3120
rect 30208 3108 30236 3139
rect 32508 3108 32536 3148
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 33505 3179 33563 3185
rect 33505 3145 33517 3179
rect 33551 3176 33563 3179
rect 34974 3176 34980 3188
rect 33551 3148 34980 3176
rect 33551 3145 33563 3148
rect 33505 3139 33563 3145
rect 34974 3136 34980 3148
rect 35032 3136 35038 3188
rect 35069 3179 35127 3185
rect 35069 3145 35081 3179
rect 35115 3176 35127 3179
rect 36722 3176 36728 3188
rect 35115 3148 36728 3176
rect 35115 3145 35127 3148
rect 35069 3139 35127 3145
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 36998 3136 37004 3188
rect 37056 3136 37062 3188
rect 30208 3080 32536 3108
rect 37090 3068 37096 3120
rect 37148 3108 37154 3120
rect 42426 3108 42432 3120
rect 37148 3080 42432 3108
rect 37148 3068 37154 3080
rect 42426 3068 42432 3080
rect 42484 3068 42490 3120
rect 54573 3111 54631 3117
rect 54573 3077 54585 3111
rect 54619 3108 54631 3111
rect 64690 3108 64696 3120
rect 54619 3080 64696 3108
rect 54619 3077 54631 3080
rect 54573 3071 54631 3077
rect 64690 3068 64696 3080
rect 64748 3068 64754 3120
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26697 3043 26755 3049
rect 26191 3012 26648 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 23014 2932 23020 2984
rect 23072 2972 23078 2984
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 23072 2944 23765 2972
rect 23072 2932 23078 2944
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 24026 2932 24032 2984
rect 24084 2972 24090 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 24084 2944 24317 2972
rect 24084 2932 24090 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 25314 2932 25320 2984
rect 25372 2932 25378 2984
rect 26234 2904 26240 2916
rect 22848 2876 26240 2904
rect 22465 2867 22523 2873
rect 26234 2864 26240 2876
rect 26292 2864 26298 2916
rect 26620 2904 26648 3012
rect 26697 3009 26709 3043
rect 26743 3009 26755 3043
rect 26697 3003 26755 3009
rect 26881 3043 26939 3049
rect 26881 3009 26893 3043
rect 26927 3040 26939 3043
rect 26970 3040 26976 3052
rect 26927 3012 26976 3040
rect 26927 3009 26939 3012
rect 26881 3003 26939 3009
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 27154 3000 27160 3052
rect 27212 3040 27218 3052
rect 27212 3012 28488 3040
rect 27212 3000 27218 3012
rect 27062 2932 27068 2984
rect 27120 2932 27126 2984
rect 27522 2932 27528 2984
rect 27580 2932 27586 2984
rect 28460 2972 28488 3012
rect 28534 3000 28540 3052
rect 28592 3000 28598 3052
rect 28644 3012 29040 3040
rect 28644 2972 28672 3012
rect 28460 2944 28672 2972
rect 28902 2932 28908 2984
rect 28960 2932 28966 2984
rect 29012 2972 29040 3012
rect 29086 3000 29092 3052
rect 29144 3000 29150 3052
rect 29546 3000 29552 3052
rect 29604 3000 29610 3052
rect 29638 3000 29644 3052
rect 29696 3040 29702 3052
rect 29733 3043 29791 3049
rect 29733 3040 29745 3043
rect 29696 3012 29745 3040
rect 29696 3000 29702 3012
rect 29733 3009 29745 3012
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 30006 3000 30012 3052
rect 30064 3000 30070 3052
rect 31478 3040 31484 3052
rect 30116 3012 31484 3040
rect 30116 2972 30144 3012
rect 31478 3000 31484 3012
rect 31536 3000 31542 3052
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 31662 3040 31668 3052
rect 31619 3012 31668 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 31662 3000 31668 3012
rect 31720 3000 31726 3052
rect 32033 3043 32091 3049
rect 32033 3009 32045 3043
rect 32079 3040 32091 3043
rect 32306 3040 32312 3052
rect 32079 3012 32312 3040
rect 32079 3009 32091 3012
rect 32033 3003 32091 3009
rect 32306 3000 32312 3012
rect 32364 3000 32370 3052
rect 32953 3043 33011 3049
rect 32953 3009 32965 3043
rect 32999 3040 33011 3043
rect 33134 3040 33140 3052
rect 32999 3012 33140 3040
rect 32999 3009 33011 3012
rect 32953 3003 33011 3009
rect 33134 3000 33140 3012
rect 33192 3000 33198 3052
rect 33318 3000 33324 3052
rect 33376 3000 33382 3052
rect 33428 3012 34008 3040
rect 29012 2944 30144 2972
rect 30190 2932 30196 2984
rect 30248 2972 30254 2984
rect 30285 2975 30343 2981
rect 30285 2972 30297 2975
rect 30248 2944 30297 2972
rect 30248 2932 30254 2944
rect 30285 2941 30297 2944
rect 30331 2941 30343 2975
rect 30285 2935 30343 2941
rect 32214 2932 32220 2984
rect 32272 2932 32278 2984
rect 29454 2904 29460 2916
rect 26620 2876 29460 2904
rect 29454 2864 29460 2876
rect 29512 2864 29518 2916
rect 29917 2907 29975 2913
rect 29917 2873 29929 2907
rect 29963 2904 29975 2907
rect 33428 2904 33456 3012
rect 33873 2975 33931 2981
rect 33873 2941 33885 2975
rect 33919 2941 33931 2975
rect 33980 2972 34008 3012
rect 34054 3000 34060 3052
rect 34112 3000 34118 3052
rect 34517 3043 34575 3049
rect 34517 3009 34529 3043
rect 34563 3040 34575 3043
rect 34606 3040 34612 3052
rect 34563 3012 34612 3040
rect 34563 3009 34575 3012
rect 34517 3003 34575 3009
rect 34606 3000 34612 3012
rect 34664 3000 34670 3052
rect 34882 3000 34888 3052
rect 34940 3000 34946 3052
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3040 35955 3043
rect 36170 3040 36176 3052
rect 35943 3012 36176 3040
rect 35943 3009 35955 3012
rect 35897 3003 35955 3009
rect 36170 3000 36176 3012
rect 36228 3000 36234 3052
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 36630 3040 36636 3052
rect 36311 3012 36636 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 36630 3000 36636 3012
rect 36688 3000 36694 3052
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 37016 3012 41414 3040
rect 34790 2972 34796 2984
rect 33980 2944 34796 2972
rect 33873 2935 33931 2941
rect 29963 2876 33456 2904
rect 33888 2904 33916 2935
rect 34790 2932 34796 2944
rect 34848 2932 34854 2984
rect 35802 2932 35808 2984
rect 35860 2932 35866 2984
rect 37016 2904 37044 3012
rect 37090 2932 37096 2984
rect 37148 2972 37154 2984
rect 41386 2972 41414 3012
rect 45922 3000 45928 3052
rect 45980 3000 45986 3052
rect 47118 3000 47124 3052
rect 47176 3040 47182 3052
rect 47489 3043 47547 3049
rect 47489 3040 47501 3043
rect 47176 3012 47501 3040
rect 47176 3000 47182 3012
rect 47489 3009 47501 3012
rect 47535 3009 47547 3043
rect 47489 3003 47547 3009
rect 49050 3000 49056 3052
rect 49108 3000 49114 3052
rect 52914 3000 52920 3052
rect 52972 3000 52978 3052
rect 53926 3000 53932 3052
rect 53984 3040 53990 3052
rect 54205 3043 54263 3049
rect 54205 3040 54217 3043
rect 53984 3012 54217 3040
rect 53984 3000 53990 3012
rect 54205 3009 54217 3012
rect 54251 3009 54263 3043
rect 54205 3003 54263 3009
rect 54662 3000 54668 3052
rect 54720 3000 54726 3052
rect 56226 3000 56232 3052
rect 56284 3000 56290 3052
rect 57790 3000 57796 3052
rect 57848 3000 57854 3052
rect 59446 3000 59452 3052
rect 59504 3000 59510 3052
rect 61194 3000 61200 3052
rect 61252 3000 61258 3052
rect 63218 3000 63224 3052
rect 63276 3000 63282 3052
rect 64782 3000 64788 3052
rect 64840 3000 64846 3052
rect 66438 3000 66444 3052
rect 66496 3000 66502 3052
rect 68094 3000 68100 3052
rect 68152 3000 68158 3052
rect 69842 3000 69848 3052
rect 69900 3000 69906 3052
rect 71406 3000 71412 3052
rect 71464 3000 71470 3052
rect 72881 3043 72939 3049
rect 72881 3009 72893 3043
rect 72927 3040 72939 3043
rect 73246 3040 73252 3052
rect 72927 3012 73252 3040
rect 72927 3009 72939 3012
rect 72881 3003 72939 3009
rect 73246 3000 73252 3012
rect 73304 3000 73310 3052
rect 63586 2972 63592 2984
rect 37148 2944 38240 2972
rect 41386 2944 63592 2972
rect 37148 2932 37154 2944
rect 33888 2876 37044 2904
rect 38212 2904 38240 2944
rect 63586 2932 63592 2944
rect 63644 2932 63650 2984
rect 44818 2904 44824 2916
rect 38212 2876 44824 2904
rect 29963 2873 29975 2876
rect 29917 2867 29975 2873
rect 44818 2864 44824 2876
rect 44876 2864 44882 2916
rect 47673 2907 47731 2913
rect 47673 2873 47685 2907
rect 47719 2904 47731 2907
rect 50062 2904 50068 2916
rect 47719 2876 50068 2904
rect 47719 2873 47731 2876
rect 47673 2867 47731 2873
rect 50062 2864 50068 2876
rect 50120 2864 50126 2916
rect 18414 2796 18420 2848
rect 18472 2796 18478 2848
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 21450 2796 21456 2848
rect 21508 2796 21514 2848
rect 22370 2796 22376 2848
rect 22428 2796 22434 2848
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 23201 2839 23259 2845
rect 23201 2836 23213 2839
rect 22612 2808 23213 2836
rect 22612 2796 22618 2808
rect 23201 2805 23213 2808
rect 23247 2805 23259 2839
rect 23201 2799 23259 2805
rect 24946 2796 24952 2848
rect 25004 2796 25010 2848
rect 25958 2796 25964 2848
rect 26016 2796 26022 2848
rect 26510 2796 26516 2848
rect 26568 2796 26574 2848
rect 28166 2796 28172 2848
rect 28224 2836 28230 2848
rect 28353 2839 28411 2845
rect 28353 2836 28365 2839
rect 28224 2808 28365 2836
rect 28224 2796 28230 2808
rect 28353 2805 28365 2808
rect 28399 2805 28411 2839
rect 28353 2799 28411 2805
rect 30926 2796 30932 2848
rect 30984 2796 30990 2848
rect 31481 2839 31539 2845
rect 31481 2805 31493 2839
rect 31527 2836 31539 2839
rect 32582 2836 32588 2848
rect 31527 2808 32588 2836
rect 31527 2805 31539 2808
rect 31481 2799 31539 2805
rect 32582 2796 32588 2808
rect 32640 2796 32646 2848
rect 32861 2839 32919 2845
rect 32861 2805 32873 2839
rect 32907 2836 32919 2839
rect 32950 2836 32956 2848
rect 32907 2808 32956 2836
rect 32907 2805 32919 2808
rect 32861 2799 32919 2805
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 33870 2796 33876 2848
rect 33928 2836 33934 2848
rect 34241 2839 34299 2845
rect 34241 2836 34253 2839
rect 33928 2808 34253 2836
rect 33928 2796 33934 2808
rect 34241 2805 34253 2808
rect 34287 2805 34299 2839
rect 34241 2799 34299 2805
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 35161 2839 35219 2845
rect 35161 2836 35173 2839
rect 34756 2808 35173 2836
rect 34756 2796 34762 2808
rect 35161 2805 35173 2808
rect 35207 2805 35219 2839
rect 35161 2799 35219 2805
rect 35802 2796 35808 2848
rect 35860 2836 35866 2848
rect 44910 2836 44916 2848
rect 35860 2808 44916 2836
rect 35860 2796 35866 2808
rect 44910 2796 44916 2808
rect 44968 2796 44974 2848
rect 46109 2839 46167 2845
rect 46109 2805 46121 2839
rect 46155 2836 46167 2839
rect 47578 2836 47584 2848
rect 46155 2808 47584 2836
rect 46155 2805 46167 2808
rect 46109 2799 46167 2805
rect 47578 2796 47584 2808
rect 47636 2796 47642 2848
rect 49237 2839 49295 2845
rect 49237 2805 49249 2839
rect 49283 2836 49295 2839
rect 52638 2836 52644 2848
rect 49283 2808 52644 2836
rect 49283 2805 49295 2808
rect 49237 2799 49295 2805
rect 52638 2796 52644 2808
rect 52696 2796 52702 2848
rect 53098 2796 53104 2848
rect 53156 2796 53162 2848
rect 54849 2839 54907 2845
rect 54849 2805 54861 2839
rect 54895 2836 54907 2839
rect 55214 2836 55220 2848
rect 54895 2808 55220 2836
rect 54895 2805 54907 2808
rect 54849 2799 54907 2805
rect 55214 2796 55220 2808
rect 55272 2796 55278 2848
rect 56410 2796 56416 2848
rect 56468 2796 56474 2848
rect 57974 2796 57980 2848
rect 58032 2796 58038 2848
rect 59633 2839 59691 2845
rect 59633 2805 59645 2839
rect 59679 2836 59691 2839
rect 60366 2836 60372 2848
rect 59679 2808 60372 2836
rect 59679 2805 59691 2808
rect 59633 2799 59691 2805
rect 60366 2796 60372 2808
rect 60424 2796 60430 2848
rect 61378 2796 61384 2848
rect 61436 2796 61442 2848
rect 63034 2796 63040 2848
rect 63092 2796 63098 2848
rect 64598 2796 64604 2848
rect 64656 2796 64662 2848
rect 66254 2796 66260 2848
rect 66312 2796 66318 2848
rect 68278 2796 68284 2848
rect 68336 2796 68342 2848
rect 69658 2796 69664 2848
rect 69716 2796 69722 2848
rect 71222 2796 71228 2848
rect 71280 2796 71286 2848
rect 73065 2839 73123 2845
rect 73065 2805 73077 2839
rect 73111 2836 73123 2839
rect 73246 2836 73252 2848
rect 73111 2808 73252 2836
rect 73111 2805 73123 2808
rect 73065 2799 73123 2805
rect 73246 2796 73252 2808
rect 73304 2796 73310 2848
rect 1012 2746 74980 2768
rect 1012 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 74980 2746
rect 1012 2672 74980 2694
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 18196 2604 18245 2632
rect 18196 2592 18202 2604
rect 18233 2601 18245 2604
rect 18279 2601 18291 2635
rect 18233 2595 18291 2601
rect 18969 2635 19027 2641
rect 18969 2601 18981 2635
rect 19015 2632 19027 2635
rect 19150 2632 19156 2644
rect 19015 2604 19156 2632
rect 19015 2601 19027 2604
rect 18969 2595 19027 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19886 2592 19892 2644
rect 19944 2592 19950 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20806 2632 20812 2644
rect 20027 2604 20812 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 21361 2635 21419 2641
rect 21361 2601 21373 2635
rect 21407 2632 21419 2635
rect 21726 2632 21732 2644
rect 21407 2604 21732 2632
rect 21407 2601 21419 2604
rect 21361 2595 21419 2601
rect 21726 2592 21732 2604
rect 21784 2592 21790 2644
rect 24026 2592 24032 2644
rect 24084 2632 24090 2644
rect 24121 2635 24179 2641
rect 24121 2632 24133 2635
rect 24084 2604 24133 2632
rect 24084 2592 24090 2604
rect 24121 2601 24133 2604
rect 24167 2601 24179 2635
rect 24121 2595 24179 2601
rect 25222 2592 25228 2644
rect 25280 2592 25286 2644
rect 25314 2592 25320 2644
rect 25372 2592 25378 2644
rect 27522 2592 27528 2644
rect 27580 2592 27586 2644
rect 29086 2592 29092 2644
rect 29144 2632 29150 2644
rect 29273 2635 29331 2641
rect 29273 2632 29285 2635
rect 29144 2604 29285 2632
rect 29144 2592 29150 2604
rect 29273 2601 29285 2604
rect 29319 2601 29331 2635
rect 70670 2632 70676 2644
rect 29273 2595 29331 2601
rect 30576 2604 70676 2632
rect 23290 2564 23296 2576
rect 17512 2536 23296 2564
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17512 2437 17540 2536
rect 23290 2524 23296 2536
rect 23348 2524 23354 2576
rect 25866 2524 25872 2576
rect 25924 2564 25930 2576
rect 30466 2564 30472 2576
rect 25924 2536 30472 2564
rect 25924 2524 25930 2536
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2496 18475 2499
rect 19702 2496 19708 2508
rect 18463 2468 19708 2496
rect 18463 2465 18475 2468
rect 18417 2459 18475 2465
rect 19702 2456 19708 2468
rect 19760 2456 19766 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 20806 2496 20812 2508
rect 20671 2468 20812 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 25958 2496 25964 2508
rect 22848 2468 25964 2496
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 17000 2400 17049 2428
rect 17000 2388 17006 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 19337 2431 19395 2437
rect 19337 2397 19349 2431
rect 19383 2428 19395 2431
rect 20162 2428 20168 2440
rect 19383 2400 20168 2428
rect 19383 2397 19395 2400
rect 19337 2391 19395 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20530 2360 20536 2372
rect 17236 2332 20536 2360
rect 17236 2301 17264 2332
rect 20530 2320 20536 2332
rect 20588 2320 20594 2372
rect 20732 2360 20760 2391
rect 21358 2388 21364 2440
rect 21416 2428 21422 2440
rect 22848 2437 22876 2468
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 27798 2456 27804 2508
rect 27856 2496 27862 2508
rect 27856 2468 28396 2496
rect 27856 2456 27862 2468
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 21416 2400 21649 2428
rect 21416 2388 21422 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 24026 2428 24032 2440
rect 23615 2400 24032 2428
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25280 2400 25881 2428
rect 25280 2388 25286 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26050 2388 26056 2440
rect 26108 2388 26114 2440
rect 26142 2388 26148 2440
rect 26200 2428 26206 2440
rect 26789 2431 26847 2437
rect 26789 2428 26801 2431
rect 26200 2400 26801 2428
rect 26200 2388 26206 2400
rect 26789 2397 26801 2400
rect 26835 2397 26847 2431
rect 26789 2391 26847 2397
rect 26878 2388 26884 2440
rect 26936 2428 26942 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26936 2400 27353 2428
rect 26936 2388 26942 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27430 2388 27436 2440
rect 27488 2428 27494 2440
rect 28368 2437 28396 2468
rect 28442 2456 28448 2508
rect 28500 2496 28506 2508
rect 30576 2496 30604 2604
rect 70670 2592 70676 2604
rect 70728 2592 70734 2644
rect 31662 2524 31668 2576
rect 31720 2524 31726 2576
rect 33134 2524 33140 2576
rect 33192 2524 33198 2576
rect 34054 2524 34060 2576
rect 34112 2564 34118 2576
rect 34241 2567 34299 2573
rect 34241 2564 34253 2567
rect 34112 2536 34253 2564
rect 34112 2524 34118 2536
rect 34241 2533 34253 2536
rect 34287 2533 34299 2567
rect 34241 2527 34299 2533
rect 34992 2536 39344 2564
rect 28500 2468 30604 2496
rect 28500 2456 28506 2468
rect 30926 2456 30932 2508
rect 30984 2456 30990 2508
rect 34992 2505 35020 2536
rect 34977 2499 35035 2505
rect 34977 2465 34989 2499
rect 35023 2465 35035 2499
rect 34977 2459 35035 2465
rect 35434 2456 35440 2508
rect 35492 2496 35498 2508
rect 36541 2499 36599 2505
rect 36541 2496 36553 2499
rect 35492 2468 36553 2496
rect 35492 2456 35498 2468
rect 36541 2465 36553 2468
rect 36587 2465 36599 2499
rect 36541 2459 36599 2465
rect 39209 2499 39267 2505
rect 39209 2465 39221 2499
rect 39255 2465 39267 2499
rect 39316 2496 39344 2536
rect 39390 2524 39396 2576
rect 39448 2564 39454 2576
rect 43346 2564 43352 2576
rect 39448 2536 43352 2564
rect 39448 2524 39454 2536
rect 43346 2524 43352 2536
rect 43404 2524 43410 2576
rect 44361 2567 44419 2573
rect 44361 2533 44373 2567
rect 44407 2564 44419 2567
rect 44726 2564 44732 2576
rect 44407 2536 44732 2564
rect 44407 2533 44419 2536
rect 44361 2527 44419 2533
rect 44726 2524 44732 2536
rect 44784 2524 44790 2576
rect 47029 2567 47087 2573
rect 47029 2533 47041 2567
rect 47075 2564 47087 2567
rect 51166 2564 51172 2576
rect 47075 2536 51172 2564
rect 47075 2533 47087 2536
rect 47029 2527 47087 2533
rect 51166 2524 51172 2536
rect 51224 2524 51230 2576
rect 53926 2524 53932 2576
rect 53984 2524 53990 2576
rect 54018 2524 54024 2576
rect 54076 2564 54082 2576
rect 63221 2567 63279 2573
rect 54076 2536 58756 2564
rect 54076 2524 54082 2536
rect 47854 2496 47860 2508
rect 39316 2468 47860 2496
rect 39209 2459 39267 2465
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 27488 2400 28089 2428
rect 27488 2388 27494 2400
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28626 2388 28632 2440
rect 28684 2388 28690 2440
rect 29178 2388 29184 2440
rect 29236 2428 29242 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29236 2400 30021 2428
rect 29236 2388 29242 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 30009 2391 30067 2397
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32490 2388 32496 2440
rect 32548 2388 32554 2440
rect 33594 2388 33600 2440
rect 33652 2388 33658 2440
rect 35161 2431 35219 2437
rect 35161 2397 35173 2431
rect 35207 2428 35219 2431
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35207 2400 35265 2428
rect 35207 2397 35219 2400
rect 35161 2391 35219 2397
rect 35253 2397 35265 2400
rect 35299 2397 35311 2431
rect 35253 2391 35311 2397
rect 35897 2431 35955 2437
rect 35897 2397 35909 2431
rect 35943 2428 35955 2431
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35943 2400 36001 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 39224 2428 39252 2459
rect 47854 2456 47860 2468
rect 47912 2456 47918 2508
rect 48038 2456 48044 2508
rect 48096 2496 48102 2508
rect 55306 2496 55312 2508
rect 48096 2468 55312 2496
rect 48096 2456 48102 2468
rect 55306 2456 55312 2468
rect 55364 2456 55370 2508
rect 55585 2499 55643 2505
rect 55585 2465 55597 2499
rect 55631 2496 55643 2499
rect 55631 2468 58664 2496
rect 55631 2465 55643 2468
rect 55585 2459 55643 2465
rect 41690 2428 41696 2440
rect 39224 2400 41696 2428
rect 35989 2391 36047 2397
rect 41690 2388 41696 2400
rect 41748 2388 41754 2440
rect 42334 2388 42340 2440
rect 42392 2428 42398 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 42392 2400 42441 2428
rect 42392 2388 42398 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 43496 2400 43729 2428
rect 43496 2388 43502 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 43717 2391 43775 2397
rect 44729 2431 44787 2437
rect 44729 2397 44741 2431
rect 44775 2428 44787 2431
rect 44913 2431 44971 2437
rect 44913 2428 44925 2431
rect 44775 2400 44925 2428
rect 44775 2397 44787 2400
rect 44729 2391 44787 2397
rect 44913 2397 44925 2400
rect 44959 2397 44971 2431
rect 44913 2391 44971 2397
rect 45554 2388 45560 2440
rect 45612 2388 45618 2440
rect 46198 2388 46204 2440
rect 46256 2388 46262 2440
rect 47302 2388 47308 2440
rect 47360 2428 47366 2440
rect 47397 2431 47455 2437
rect 47397 2428 47409 2431
rect 47360 2400 47409 2428
rect 47360 2388 47366 2400
rect 47397 2397 47409 2400
rect 47443 2397 47455 2431
rect 47397 2391 47455 2397
rect 47780 2400 48084 2428
rect 21726 2360 21732 2372
rect 20732 2332 21732 2360
rect 21726 2320 21732 2332
rect 21784 2320 21790 2372
rect 23201 2363 23259 2369
rect 23201 2329 23213 2363
rect 23247 2360 23259 2363
rect 23247 2332 36584 2360
rect 23247 2329 23259 2332
rect 23201 2323 23259 2329
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17313 2295 17371 2301
rect 17313 2261 17325 2295
rect 17359 2292 17371 2295
rect 17770 2292 17776 2304
rect 17359 2264 17776 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 20898 2292 20904 2304
rect 17920 2264 20904 2292
rect 17920 2252 17926 2264
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 26694 2252 26700 2304
rect 26752 2252 26758 2304
rect 28534 2252 28540 2304
rect 28592 2252 28598 2304
rect 29086 2252 29092 2304
rect 29144 2292 29150 2304
rect 29457 2295 29515 2301
rect 29457 2292 29469 2295
rect 29144 2264 29469 2292
rect 29144 2252 29150 2264
rect 29457 2261 29469 2264
rect 29503 2261 29515 2295
rect 29457 2255 29515 2261
rect 30282 2252 30288 2304
rect 30340 2252 30346 2304
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 31757 2295 31815 2301
rect 31757 2292 31769 2295
rect 31352 2264 31769 2292
rect 31352 2252 31358 2264
rect 31757 2261 31769 2264
rect 31803 2261 31815 2295
rect 31757 2255 31815 2261
rect 33042 2252 33048 2304
rect 33100 2292 33106 2304
rect 35066 2292 35072 2304
rect 33100 2264 35072 2292
rect 33100 2252 33106 2264
rect 35066 2252 35072 2264
rect 35124 2252 35130 2304
rect 36556 2292 36584 2332
rect 39114 2320 39120 2372
rect 39172 2360 39178 2372
rect 39485 2363 39543 2369
rect 39485 2360 39497 2363
rect 39172 2332 39497 2360
rect 39172 2320 39178 2332
rect 39485 2329 39497 2332
rect 39531 2329 39543 2363
rect 39485 2323 39543 2329
rect 43070 2320 43076 2372
rect 43128 2320 43134 2372
rect 46382 2360 46388 2372
rect 43180 2332 46388 2360
rect 39390 2292 39396 2304
rect 36556 2264 39396 2292
rect 39390 2252 39396 2264
rect 39448 2252 39454 2304
rect 39574 2252 39580 2304
rect 39632 2292 39638 2304
rect 43180 2292 43208 2332
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 46676 2332 46980 2360
rect 39632 2264 43208 2292
rect 44545 2295 44603 2301
rect 39632 2252 39638 2264
rect 44545 2261 44557 2295
rect 44591 2292 44603 2295
rect 46676 2292 46704 2332
rect 44591 2264 46704 2292
rect 46753 2295 46811 2301
rect 44591 2261 44603 2264
rect 44545 2255 44603 2261
rect 46753 2261 46765 2295
rect 46799 2292 46811 2295
rect 46842 2292 46848 2304
rect 46799 2264 46848 2292
rect 46799 2261 46811 2264
rect 46753 2255 46811 2261
rect 46842 2252 46848 2264
rect 46900 2252 46906 2304
rect 46952 2292 46980 2332
rect 47210 2320 47216 2372
rect 47268 2320 47274 2372
rect 47780 2292 47808 2400
rect 48056 2360 48084 2400
rect 49050 2388 49056 2440
rect 49108 2388 49114 2440
rect 53377 2431 53435 2437
rect 53377 2397 53389 2431
rect 53423 2428 53435 2431
rect 53834 2428 53840 2440
rect 53423 2400 53840 2428
rect 53423 2397 53435 2400
rect 53377 2391 53435 2397
rect 53834 2388 53840 2400
rect 53892 2388 53898 2440
rect 53926 2388 53932 2440
rect 53984 2428 53990 2440
rect 54113 2431 54171 2437
rect 54113 2428 54125 2431
rect 53984 2400 54125 2428
rect 53984 2388 53990 2400
rect 54113 2397 54125 2400
rect 54159 2397 54171 2431
rect 54113 2391 54171 2397
rect 57330 2388 57336 2440
rect 57388 2388 57394 2440
rect 53742 2360 53748 2372
rect 48056 2332 53748 2360
rect 53742 2320 53748 2332
rect 53800 2320 53806 2372
rect 55030 2320 55036 2372
rect 55088 2360 55094 2372
rect 55309 2363 55367 2369
rect 55309 2360 55321 2363
rect 55088 2332 55321 2360
rect 55088 2320 55094 2332
rect 55309 2329 55321 2332
rect 55355 2329 55367 2363
rect 55309 2323 55367 2329
rect 56137 2363 56195 2369
rect 56137 2329 56149 2363
rect 56183 2360 56195 2363
rect 56686 2360 56692 2372
rect 56183 2332 56692 2360
rect 56183 2329 56195 2332
rect 56137 2323 56195 2329
rect 56686 2320 56692 2332
rect 56744 2320 56750 2372
rect 58636 2360 58664 2468
rect 58728 2428 58756 2536
rect 63221 2533 63233 2567
rect 63267 2564 63279 2567
rect 66162 2564 66168 2576
rect 63267 2536 66168 2564
rect 63267 2533 63279 2536
rect 63221 2527 63279 2533
rect 66162 2524 66168 2536
rect 66220 2524 66226 2576
rect 60737 2499 60795 2505
rect 60737 2465 60749 2499
rect 60783 2496 60795 2499
rect 65702 2496 65708 2508
rect 60783 2468 65708 2496
rect 60783 2465 60795 2468
rect 60737 2459 60795 2465
rect 65702 2456 65708 2468
rect 65760 2456 65766 2508
rect 67450 2456 67456 2508
rect 67508 2456 67514 2508
rect 58728 2400 61148 2428
rect 60734 2360 60740 2372
rect 57808 2332 58572 2360
rect 58636 2332 60740 2360
rect 46952 2264 47808 2292
rect 48041 2295 48099 2301
rect 48041 2261 48053 2295
rect 48087 2292 48099 2295
rect 49418 2292 49424 2304
rect 48087 2264 49424 2292
rect 48087 2261 48099 2264
rect 48041 2255 48099 2261
rect 49418 2252 49424 2264
rect 49476 2252 49482 2304
rect 49510 2252 49516 2304
rect 49568 2292 49574 2304
rect 49697 2295 49755 2301
rect 49697 2292 49709 2295
rect 49568 2264 49709 2292
rect 49568 2252 49574 2264
rect 49697 2261 49709 2264
rect 49743 2261 49755 2295
rect 49697 2255 49755 2261
rect 54754 2252 54760 2304
rect 54812 2252 54818 2304
rect 56045 2295 56103 2301
rect 56045 2261 56057 2295
rect 56091 2292 56103 2295
rect 57808 2292 57836 2332
rect 56091 2264 57836 2292
rect 56091 2261 56103 2264
rect 56045 2255 56103 2261
rect 57882 2252 57888 2304
rect 57940 2292 57946 2304
rect 57977 2295 58035 2301
rect 57977 2292 57989 2295
rect 57940 2264 57989 2292
rect 57940 2252 57946 2264
rect 57977 2261 57989 2264
rect 58023 2261 58035 2295
rect 58544 2292 58572 2332
rect 60734 2320 60740 2332
rect 60792 2320 60798 2372
rect 61010 2320 61016 2372
rect 61068 2320 61074 2372
rect 61120 2360 61148 2400
rect 62298 2388 62304 2440
rect 62356 2388 62362 2440
rect 62408 2400 64874 2428
rect 62408 2360 62436 2400
rect 63405 2363 63463 2369
rect 61120 2332 62436 2360
rect 62868 2332 63356 2360
rect 62868 2292 62896 2332
rect 58544 2264 62896 2292
rect 57977 2255 58035 2261
rect 62942 2252 62948 2304
rect 63000 2252 63006 2304
rect 63328 2292 63356 2332
rect 63405 2329 63417 2363
rect 63451 2360 63463 2363
rect 63586 2360 63592 2372
rect 63451 2332 63592 2360
rect 63451 2329 63463 2332
rect 63405 2323 63463 2329
rect 63586 2320 63592 2332
rect 63644 2320 63650 2372
rect 64846 2360 64874 2400
rect 65518 2388 65524 2440
rect 65576 2428 65582 2440
rect 65613 2431 65671 2437
rect 65613 2428 65625 2431
rect 65576 2400 65625 2428
rect 65576 2388 65582 2400
rect 65613 2397 65625 2400
rect 65659 2397 65671 2431
rect 65613 2391 65671 2397
rect 67266 2388 67272 2440
rect 67324 2428 67330 2440
rect 67729 2431 67787 2437
rect 67729 2428 67741 2431
rect 67324 2400 67741 2428
rect 67324 2388 67330 2400
rect 67729 2397 67741 2400
rect 67775 2397 67787 2431
rect 67729 2391 67787 2397
rect 69934 2388 69940 2440
rect 69992 2388 69998 2440
rect 70486 2388 70492 2440
rect 70544 2428 70550 2440
rect 70673 2431 70731 2437
rect 70673 2428 70685 2431
rect 70544 2400 70685 2428
rect 70544 2388 70550 2400
rect 70673 2397 70685 2400
rect 70719 2397 70731 2431
rect 70673 2391 70731 2397
rect 67542 2360 67548 2372
rect 64846 2332 67548 2360
rect 67542 2320 67548 2332
rect 67600 2320 67606 2372
rect 63678 2292 63684 2304
rect 63328 2264 63684 2292
rect 63678 2252 63684 2264
rect 63736 2252 63742 2304
rect 66070 2252 66076 2304
rect 66128 2292 66134 2304
rect 66257 2295 66315 2301
rect 66257 2292 66269 2295
rect 66128 2264 66269 2292
rect 66128 2252 66134 2264
rect 66257 2261 66269 2264
rect 66303 2261 66315 2295
rect 66257 2255 66315 2261
rect 69293 2295 69351 2301
rect 69293 2261 69305 2295
rect 69339 2292 69351 2295
rect 69382 2292 69388 2304
rect 69339 2264 69388 2292
rect 69339 2261 69351 2264
rect 69293 2255 69351 2261
rect 69382 2252 69388 2264
rect 69440 2252 69446 2304
rect 71038 2252 71044 2304
rect 71096 2292 71102 2304
rect 71317 2295 71375 2301
rect 71317 2292 71329 2295
rect 71096 2264 71329 2292
rect 71096 2252 71102 2264
rect 71317 2261 71329 2264
rect 71363 2261 71375 2295
rect 71317 2255 71375 2261
rect 1012 2202 74980 2224
rect 1012 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74980 2202
rect 1012 2128 74980 2150
rect 16393 2091 16451 2097
rect 16393 2057 16405 2091
rect 16439 2057 16451 2091
rect 16393 2051 16451 2057
rect 17405 2091 17463 2097
rect 17405 2057 17417 2091
rect 17451 2088 17463 2091
rect 17586 2088 17592 2100
rect 17451 2060 17592 2088
rect 17451 2057 17463 2060
rect 17405 2051 17463 2057
rect 16408 2020 16436 2051
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 18141 2091 18199 2097
rect 18141 2057 18153 2091
rect 18187 2088 18199 2091
rect 18230 2088 18236 2100
rect 18187 2060 18236 2088
rect 18187 2057 18199 2060
rect 18141 2051 18199 2057
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 21450 2088 21456 2100
rect 19904 2060 21456 2088
rect 17862 2020 17868 2032
rect 16408 1992 17868 2020
rect 17862 1980 17868 1992
rect 17920 1980 17926 2032
rect 19904 2020 19932 2060
rect 21450 2048 21456 2060
rect 21508 2048 21514 2100
rect 24121 2091 24179 2097
rect 24121 2057 24133 2091
rect 24167 2088 24179 2091
rect 24578 2088 24584 2100
rect 24167 2060 24584 2088
rect 24167 2057 24179 2060
rect 24121 2051 24179 2057
rect 24578 2048 24584 2060
rect 24636 2048 24642 2100
rect 31849 2091 31907 2097
rect 28092 2060 31754 2088
rect 28092 2029 28120 2060
rect 28077 2023 28135 2029
rect 19274 1992 19932 2020
rect 19996 1992 27016 2020
rect 16209 1955 16267 1961
rect 16209 1921 16221 1955
rect 16255 1952 16267 1955
rect 16390 1952 16396 1964
rect 16255 1924 16396 1952
rect 16255 1921 16267 1924
rect 16209 1915 16267 1921
rect 16390 1912 16396 1924
rect 16448 1912 16454 1964
rect 17589 1955 17647 1961
rect 17589 1921 17601 1955
rect 17635 1952 17647 1955
rect 18414 1952 18420 1964
rect 17635 1924 18420 1952
rect 17635 1921 17647 1924
rect 17589 1915 17647 1921
rect 18414 1912 18420 1924
rect 18472 1912 18478 1964
rect 19996 1961 20024 1992
rect 19981 1955 20039 1961
rect 19981 1921 19993 1955
rect 20027 1921 20039 1955
rect 19981 1915 20039 1921
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 21450 1912 21456 1964
rect 21508 1912 21514 1964
rect 22189 1955 22247 1961
rect 21560 1924 21772 1952
rect 16853 1887 16911 1893
rect 16853 1853 16865 1887
rect 16899 1884 16911 1887
rect 18046 1884 18052 1896
rect 16899 1856 18052 1884
rect 16899 1853 16911 1856
rect 16853 1847 16911 1853
rect 18046 1844 18052 1856
rect 18104 1844 18110 1896
rect 19705 1887 19763 1893
rect 19705 1853 19717 1887
rect 19751 1884 19763 1887
rect 21560 1884 21588 1924
rect 19751 1856 21588 1884
rect 21744 1884 21772 1924
rect 22189 1921 22201 1955
rect 22235 1952 22247 1955
rect 22370 1952 22376 1964
rect 22235 1924 22376 1952
rect 22235 1921 22247 1924
rect 22189 1915 22247 1921
rect 22370 1912 22376 1924
rect 22428 1912 22434 1964
rect 23474 1952 23480 1964
rect 22756 1924 23480 1952
rect 22756 1884 22784 1924
rect 23474 1912 23480 1924
rect 23532 1912 23538 1964
rect 24397 1955 24455 1961
rect 24397 1921 24409 1955
rect 24443 1952 24455 1955
rect 24946 1952 24952 1964
rect 24443 1924 24952 1952
rect 24443 1921 24455 1924
rect 24397 1915 24455 1921
rect 24946 1912 24952 1924
rect 25004 1912 25010 1964
rect 25866 1912 25872 1964
rect 25924 1912 25930 1964
rect 26142 1912 26148 1964
rect 26200 1912 26206 1964
rect 26694 1912 26700 1964
rect 26752 1952 26758 1964
rect 26881 1955 26939 1961
rect 26881 1952 26893 1955
rect 26752 1924 26893 1952
rect 26752 1912 26758 1924
rect 26881 1921 26893 1924
rect 26927 1921 26939 1955
rect 26988 1952 27016 1992
rect 28077 1989 28089 2023
rect 28123 1989 28135 2023
rect 28077 1983 28135 1989
rect 28534 1980 28540 2032
rect 28592 2020 28598 2032
rect 31726 2020 31754 2060
rect 31849 2057 31861 2091
rect 31895 2088 31907 2091
rect 32306 2088 32312 2100
rect 31895 2060 32312 2088
rect 31895 2057 31907 2060
rect 31849 2051 31907 2057
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 32490 2048 32496 2100
rect 32548 2048 32554 2100
rect 34606 2048 34612 2100
rect 34664 2048 34670 2100
rect 36630 2048 36636 2100
rect 36688 2088 36694 2100
rect 36817 2091 36875 2097
rect 36817 2088 36829 2091
rect 36688 2060 36829 2088
rect 36688 2048 36694 2060
rect 36817 2057 36829 2060
rect 36863 2057 36875 2091
rect 36817 2051 36875 2057
rect 39114 2048 39120 2100
rect 39172 2048 39178 2100
rect 41690 2048 41696 2100
rect 41748 2088 41754 2100
rect 47026 2088 47032 2100
rect 41748 2060 47032 2088
rect 41748 2048 41754 2060
rect 47026 2048 47032 2060
rect 47084 2048 47090 2100
rect 47121 2091 47179 2097
rect 47121 2057 47133 2091
rect 47167 2088 47179 2091
rect 48038 2088 48044 2100
rect 47167 2060 48044 2088
rect 47167 2057 47179 2060
rect 47121 2051 47179 2057
rect 48038 2048 48044 2060
rect 48096 2048 48102 2100
rect 52273 2091 52331 2097
rect 52273 2057 52285 2091
rect 52319 2088 52331 2091
rect 54018 2088 54024 2100
rect 52319 2060 54024 2088
rect 52319 2057 52331 2060
rect 52273 2051 52331 2057
rect 54018 2048 54024 2060
rect 54076 2048 54082 2100
rect 55030 2048 55036 2100
rect 55088 2048 55094 2100
rect 58897 2091 58955 2097
rect 58897 2057 58909 2091
rect 58943 2088 58955 2091
rect 61470 2088 61476 2100
rect 58943 2060 61476 2088
rect 58943 2057 58955 2060
rect 58897 2051 58955 2057
rect 61470 2048 61476 2060
rect 61528 2048 61534 2100
rect 63586 2048 63592 2100
rect 63644 2048 63650 2100
rect 64846 2060 67128 2088
rect 64846 2020 64874 2060
rect 28592 1992 29776 2020
rect 31726 1992 64874 2020
rect 28592 1980 28598 1992
rect 28905 1955 28963 1961
rect 26988 1924 28856 1952
rect 26881 1915 26939 1921
rect 21744 1856 22784 1884
rect 19751 1853 19763 1856
rect 19705 1847 19763 1853
rect 22830 1844 22836 1896
rect 22888 1844 22894 1896
rect 23569 1887 23627 1893
rect 23569 1853 23581 1887
rect 23615 1884 23627 1887
rect 24670 1884 24676 1896
rect 23615 1856 24676 1884
rect 23615 1853 23627 1856
rect 23569 1847 23627 1853
rect 24670 1844 24676 1856
rect 24728 1844 24734 1896
rect 25409 1887 25467 1893
rect 25409 1853 25421 1887
rect 25455 1884 25467 1887
rect 28442 1884 28448 1896
rect 25455 1856 28448 1884
rect 25455 1853 25467 1856
rect 25409 1847 25467 1853
rect 28442 1844 28448 1856
rect 28500 1844 28506 1896
rect 28721 1887 28779 1893
rect 28721 1853 28733 1887
rect 28767 1853 28779 1887
rect 28721 1847 28779 1853
rect 21450 1776 21456 1828
rect 21508 1816 21514 1828
rect 25685 1819 25743 1825
rect 25685 1816 25697 1819
rect 21508 1788 25697 1816
rect 21508 1776 21514 1788
rect 25685 1785 25697 1788
rect 25731 1785 25743 1819
rect 25685 1779 25743 1785
rect 18233 1751 18291 1757
rect 18233 1717 18245 1751
rect 18279 1748 18291 1751
rect 20622 1748 20628 1760
rect 18279 1720 20628 1748
rect 18279 1717 18291 1720
rect 18233 1711 18291 1717
rect 20622 1708 20628 1720
rect 20680 1708 20686 1760
rect 26697 1751 26755 1757
rect 26697 1717 26709 1751
rect 26743 1748 26755 1751
rect 26970 1748 26976 1760
rect 26743 1720 26976 1748
rect 26743 1717 26755 1720
rect 26697 1711 26755 1717
rect 26970 1708 26976 1720
rect 27028 1708 27034 1760
rect 28736 1748 28764 1847
rect 28828 1816 28856 1924
rect 28905 1921 28917 1955
rect 28951 1921 28963 1955
rect 28905 1915 28963 1921
rect 28920 1884 28948 1915
rect 29086 1912 29092 1964
rect 29144 1912 29150 1964
rect 29546 1912 29552 1964
rect 29604 1952 29610 1964
rect 29748 1961 29776 1992
rect 66898 1980 66904 2032
rect 66956 2020 66962 2032
rect 66993 2023 67051 2029
rect 66993 2020 67005 2023
rect 66956 1992 67005 2020
rect 66956 1980 66962 1992
rect 66993 1989 67005 1992
rect 67039 1989 67051 2023
rect 67100 2020 67128 2060
rect 67266 2048 67272 2100
rect 67324 2048 67330 2100
rect 70578 2088 70584 2100
rect 67744 2060 70584 2088
rect 67744 2020 67772 2060
rect 70578 2048 70584 2060
rect 70636 2048 70642 2100
rect 67100 1992 67772 2020
rect 69109 2023 69167 2029
rect 66993 1983 67051 1989
rect 69109 1989 69121 2023
rect 69155 2020 69167 2023
rect 69198 2020 69204 2032
rect 69155 1992 69204 2020
rect 69155 1989 69167 1992
rect 69109 1983 69167 1989
rect 69198 1980 69204 1992
rect 69256 1980 69262 2032
rect 70118 1980 70124 2032
rect 70176 2020 70182 2032
rect 71961 2023 72019 2029
rect 71961 2020 71973 2023
rect 70176 1992 71973 2020
rect 70176 1980 70182 1992
rect 71961 1989 71973 1992
rect 72007 1989 72019 2023
rect 71961 1983 72019 1989
rect 29641 1955 29699 1961
rect 29641 1952 29653 1955
rect 29604 1924 29653 1952
rect 29604 1912 29610 1924
rect 29641 1921 29653 1924
rect 29687 1921 29699 1955
rect 29641 1915 29699 1921
rect 29733 1955 29791 1961
rect 29733 1921 29745 1955
rect 29779 1921 29791 1955
rect 29733 1915 29791 1921
rect 29914 1912 29920 1964
rect 29972 1952 29978 1964
rect 29972 1924 30420 1952
rect 29972 1912 29978 1924
rect 30282 1884 30288 1896
rect 28920 1856 30288 1884
rect 30282 1844 30288 1856
rect 30340 1844 30346 1896
rect 30392 1893 30420 1924
rect 31294 1912 31300 1964
rect 31352 1912 31358 1964
rect 33321 1955 33379 1961
rect 33321 1921 33333 1955
rect 33367 1952 33379 1955
rect 34054 1952 34060 1964
rect 33367 1924 34060 1952
rect 33367 1921 33379 1924
rect 33321 1915 33379 1921
rect 34054 1912 34060 1924
rect 34112 1912 34118 1964
rect 34790 1912 34796 1964
rect 34848 1912 34854 1964
rect 38105 1955 38163 1961
rect 38105 1921 38117 1955
rect 38151 1952 38163 1955
rect 38289 1955 38347 1961
rect 38289 1952 38301 1955
rect 38151 1924 38301 1952
rect 38151 1921 38163 1924
rect 38105 1915 38163 1921
rect 38289 1921 38301 1924
rect 38335 1921 38347 1955
rect 38289 1915 38347 1921
rect 39022 1912 39028 1964
rect 39080 1952 39086 1964
rect 40405 1955 40463 1961
rect 40405 1952 40417 1955
rect 39080 1924 40417 1952
rect 39080 1912 39086 1924
rect 40405 1921 40417 1924
rect 40451 1921 40463 1955
rect 40405 1915 40463 1921
rect 41693 1955 41751 1961
rect 41693 1921 41705 1955
rect 41739 1952 41751 1955
rect 41785 1955 41843 1961
rect 41785 1952 41797 1955
rect 41739 1924 41797 1952
rect 41739 1921 41751 1924
rect 41693 1915 41751 1921
rect 41785 1921 41797 1924
rect 41831 1921 41843 1955
rect 41785 1915 41843 1921
rect 42705 1955 42763 1961
rect 42705 1921 42717 1955
rect 42751 1952 42763 1955
rect 42886 1952 42892 1964
rect 42751 1924 42892 1952
rect 42751 1921 42763 1924
rect 42705 1915 42763 1921
rect 42886 1912 42892 1924
rect 42944 1912 42950 1964
rect 42978 1912 42984 1964
rect 43036 1912 43042 1964
rect 44729 1955 44787 1961
rect 43364 1924 43576 1952
rect 30377 1887 30435 1893
rect 30377 1853 30389 1887
rect 30423 1853 30435 1887
rect 30377 1847 30435 1853
rect 32398 1844 32404 1896
rect 32456 1884 32462 1896
rect 33137 1887 33195 1893
rect 33137 1884 33149 1887
rect 32456 1856 33149 1884
rect 32456 1844 32462 1856
rect 33137 1853 33149 1856
rect 33183 1853 33195 1887
rect 33137 1847 33195 1853
rect 33873 1887 33931 1893
rect 33873 1853 33885 1887
rect 33919 1884 33931 1887
rect 33965 1887 34023 1893
rect 33965 1884 33977 1887
rect 33919 1856 33977 1884
rect 33919 1853 33931 1856
rect 33873 1847 33931 1853
rect 33965 1853 33977 1856
rect 34011 1853 34023 1887
rect 33965 1847 34023 1853
rect 34606 1844 34612 1896
rect 34664 1884 34670 1896
rect 35161 1887 35219 1893
rect 35161 1884 35173 1887
rect 34664 1856 35173 1884
rect 34664 1844 34670 1856
rect 35161 1853 35173 1856
rect 35207 1853 35219 1887
rect 35161 1847 35219 1853
rect 36170 1844 36176 1896
rect 36228 1844 36234 1896
rect 37550 1844 37556 1896
rect 37608 1844 37614 1896
rect 39761 1887 39819 1893
rect 39761 1853 39773 1887
rect 39807 1884 39819 1887
rect 39853 1887 39911 1893
rect 39853 1884 39865 1887
rect 39807 1856 39865 1884
rect 39807 1853 39819 1856
rect 39761 1847 39819 1853
rect 39853 1853 39865 1856
rect 39899 1853 39911 1887
rect 39853 1847 39911 1853
rect 41138 1844 41144 1896
rect 41196 1844 41202 1896
rect 43364 1884 43392 1924
rect 42904 1856 43392 1884
rect 43441 1887 43499 1893
rect 35894 1816 35900 1828
rect 28828 1788 35900 1816
rect 35894 1776 35900 1788
rect 35952 1776 35958 1828
rect 38565 1819 38623 1825
rect 38565 1785 38577 1819
rect 38611 1816 38623 1819
rect 42904 1816 42932 1856
rect 43441 1853 43453 1887
rect 43487 1853 43499 1887
rect 43441 1847 43499 1853
rect 38611 1788 42932 1816
rect 38611 1785 38623 1788
rect 38565 1779 38623 1785
rect 42978 1776 42984 1828
rect 43036 1816 43042 1828
rect 43456 1816 43484 1847
rect 43036 1788 43484 1816
rect 43548 1816 43576 1924
rect 44729 1921 44741 1955
rect 44775 1952 44787 1955
rect 44775 1924 45048 1952
rect 44775 1921 44787 1924
rect 44729 1915 44787 1921
rect 44910 1844 44916 1896
rect 44968 1844 44974 1896
rect 45020 1884 45048 1924
rect 45370 1912 45376 1964
rect 45428 1912 45434 1964
rect 45646 1912 45652 1964
rect 45704 1952 45710 1964
rect 46753 1955 46811 1961
rect 46753 1952 46765 1955
rect 45704 1924 46765 1952
rect 45704 1912 45710 1924
rect 46753 1921 46765 1924
rect 46799 1921 46811 1955
rect 46753 1915 46811 1921
rect 46842 1912 46848 1964
rect 46900 1952 46906 1964
rect 46937 1955 46995 1961
rect 46937 1952 46949 1955
rect 46900 1924 46949 1952
rect 46900 1912 46906 1924
rect 46937 1921 46949 1924
rect 46983 1921 46995 1955
rect 46937 1915 46995 1921
rect 47578 1912 47584 1964
rect 47636 1952 47642 1964
rect 47949 1955 48007 1961
rect 47949 1952 47961 1955
rect 47636 1924 47961 1952
rect 47636 1912 47642 1924
rect 47949 1921 47961 1924
rect 47995 1921 48007 1955
rect 47949 1915 48007 1921
rect 49510 1912 49516 1964
rect 49568 1912 49574 1964
rect 50065 1955 50123 1961
rect 50065 1921 50077 1955
rect 50111 1952 50123 1955
rect 50249 1955 50307 1961
rect 50249 1952 50261 1955
rect 50111 1924 50261 1952
rect 50111 1921 50123 1924
rect 50065 1915 50123 1921
rect 50249 1921 50261 1924
rect 50295 1921 50307 1955
rect 50249 1915 50307 1921
rect 51813 1955 51871 1961
rect 51813 1921 51825 1955
rect 51859 1952 51871 1955
rect 51997 1955 52055 1961
rect 51997 1952 52009 1955
rect 51859 1924 52009 1952
rect 51859 1921 51871 1924
rect 51813 1915 51871 1921
rect 51997 1921 52009 1924
rect 52043 1921 52055 1955
rect 51997 1915 52055 1921
rect 53098 1912 53104 1964
rect 53156 1912 53162 1964
rect 54481 1955 54539 1961
rect 54481 1921 54493 1955
rect 54527 1952 54539 1955
rect 54754 1952 54760 1964
rect 54527 1924 54760 1952
rect 54527 1921 54539 1924
rect 54481 1915 54539 1921
rect 54754 1912 54760 1924
rect 54812 1912 54818 1964
rect 56410 1912 56416 1964
rect 56468 1912 56474 1964
rect 57882 1912 57888 1964
rect 57940 1912 57946 1964
rect 58437 1955 58495 1961
rect 58437 1921 58449 1955
rect 58483 1952 58495 1955
rect 58621 1955 58679 1961
rect 58621 1952 58633 1955
rect 58483 1924 58633 1952
rect 58483 1921 58495 1924
rect 58437 1915 58495 1921
rect 58621 1921 58633 1924
rect 58667 1921 58679 1955
rect 58621 1915 58679 1921
rect 59817 1955 59875 1961
rect 59817 1921 59829 1955
rect 59863 1952 59875 1955
rect 60001 1955 60059 1961
rect 60001 1952 60013 1955
rect 59863 1924 60013 1952
rect 59863 1921 59875 1924
rect 59817 1915 59875 1921
rect 60001 1921 60013 1924
rect 60047 1921 60059 1955
rect 60001 1915 60059 1921
rect 61378 1912 61384 1964
rect 61436 1912 61442 1964
rect 62942 1912 62948 1964
rect 63000 1912 63006 1964
rect 64598 1912 64604 1964
rect 64656 1912 64662 1964
rect 66070 1912 66076 1964
rect 66128 1912 66134 1964
rect 66625 1955 66683 1961
rect 66625 1921 66637 1955
rect 66671 1952 66683 1955
rect 66717 1955 66775 1961
rect 66717 1952 66729 1955
rect 66671 1924 66729 1952
rect 66671 1921 66683 1924
rect 66625 1915 66683 1921
rect 66717 1921 66729 1924
rect 66763 1921 66775 1955
rect 66717 1915 66775 1921
rect 67174 1912 67180 1964
rect 67232 1952 67238 1964
rect 68649 1955 68707 1961
rect 68649 1952 68661 1955
rect 67232 1924 68661 1952
rect 67232 1912 67238 1924
rect 68649 1921 68661 1924
rect 68695 1921 68707 1955
rect 68649 1915 68707 1921
rect 69382 1912 69388 1964
rect 69440 1912 69446 1964
rect 69658 1912 69664 1964
rect 69716 1912 69722 1964
rect 71038 1912 71044 1964
rect 71096 1912 71102 1964
rect 71593 1955 71651 1961
rect 71593 1921 71605 1955
rect 71639 1952 71651 1955
rect 71685 1955 71743 1961
rect 71685 1952 71697 1955
rect 71639 1924 71697 1952
rect 71639 1921 71651 1924
rect 71593 1915 71651 1921
rect 71685 1921 71697 1924
rect 71731 1921 71743 1955
rect 71685 1915 71743 1921
rect 45465 1887 45523 1893
rect 45465 1884 45477 1887
rect 45020 1856 45477 1884
rect 45465 1853 45477 1856
rect 45511 1853 45523 1887
rect 45465 1847 45523 1853
rect 46014 1844 46020 1896
rect 46072 1844 46078 1896
rect 46198 1844 46204 1896
rect 46256 1844 46262 1896
rect 47854 1844 47860 1896
rect 47912 1884 47918 1896
rect 48409 1887 48467 1893
rect 48409 1884 48421 1887
rect 47912 1856 48421 1884
rect 47912 1844 47918 1856
rect 48409 1853 48421 1856
rect 48455 1853 48467 1887
rect 48409 1847 48467 1853
rect 51258 1844 51264 1896
rect 51316 1844 51322 1896
rect 51828 1856 52868 1884
rect 50430 1816 50436 1828
rect 43548 1788 50436 1816
rect 43036 1776 43042 1788
rect 50430 1776 50436 1788
rect 50488 1776 50494 1828
rect 50525 1819 50583 1825
rect 50525 1785 50537 1819
rect 50571 1816 50583 1819
rect 51828 1816 51856 1856
rect 52730 1816 52736 1828
rect 50571 1788 51856 1816
rect 51920 1788 52736 1816
rect 50571 1785 50583 1788
rect 50525 1779 50583 1785
rect 39574 1748 39580 1760
rect 28736 1720 39580 1748
rect 39574 1708 39580 1720
rect 39632 1708 39638 1760
rect 41969 1751 42027 1757
rect 41969 1717 41981 1751
rect 42015 1748 42027 1751
rect 42242 1748 42248 1760
rect 42015 1720 42248 1748
rect 42015 1717 42027 1720
rect 41969 1711 42027 1717
rect 42242 1708 42248 1720
rect 42300 1708 42306 1760
rect 42521 1751 42579 1757
rect 42521 1717 42533 1751
rect 42567 1748 42579 1751
rect 51920 1748 51948 1788
rect 52730 1776 52736 1788
rect 52788 1776 52794 1828
rect 52840 1816 52868 1856
rect 52914 1844 52920 1896
rect 52972 1884 52978 1896
rect 53377 1887 53435 1893
rect 53377 1884 53389 1887
rect 52972 1856 53389 1884
rect 52972 1844 52978 1856
rect 53377 1853 53389 1856
rect 53423 1853 53435 1887
rect 53377 1847 53435 1853
rect 55582 1844 55588 1896
rect 55640 1844 55646 1896
rect 56134 1844 56140 1896
rect 56192 1884 56198 1896
rect 56689 1887 56747 1893
rect 56689 1884 56701 1887
rect 56192 1856 56701 1884
rect 56192 1844 56198 1856
rect 56689 1853 56701 1856
rect 56735 1853 56747 1887
rect 56689 1847 56747 1853
rect 59265 1887 59323 1893
rect 59265 1853 59277 1887
rect 59311 1884 59323 1887
rect 59354 1884 59360 1896
rect 59311 1856 59360 1884
rect 59311 1853 59323 1856
rect 59265 1847 59323 1853
rect 59354 1844 59360 1856
rect 59412 1844 59418 1896
rect 60550 1844 60556 1896
rect 60608 1844 60614 1896
rect 61102 1844 61108 1896
rect 61160 1884 61166 1896
rect 61657 1887 61715 1893
rect 61657 1884 61669 1887
rect 61160 1856 61669 1884
rect 61160 1844 61166 1856
rect 61657 1853 61669 1856
rect 61703 1853 61715 1887
rect 61657 1847 61715 1853
rect 63862 1844 63868 1896
rect 63920 1844 63926 1896
rect 64690 1844 64696 1896
rect 64748 1884 64754 1896
rect 64969 1887 65027 1893
rect 64969 1884 64981 1887
rect 64748 1856 64981 1884
rect 64748 1844 64754 1856
rect 64969 1853 64981 1856
rect 65015 1853 65027 1887
rect 64969 1847 65027 1853
rect 67913 1887 67971 1893
rect 67913 1853 67925 1887
rect 67959 1884 67971 1887
rect 68097 1887 68155 1893
rect 68097 1884 68109 1887
rect 67959 1856 68109 1884
rect 67959 1853 67971 1856
rect 67913 1847 67971 1853
rect 68097 1853 68109 1856
rect 68143 1853 68155 1887
rect 69937 1887 69995 1893
rect 69937 1884 69949 1887
rect 68097 1847 68155 1853
rect 69400 1856 69949 1884
rect 69400 1828 69428 1856
rect 69937 1853 69949 1856
rect 69983 1853 69995 1887
rect 69937 1847 69995 1853
rect 72234 1844 72240 1896
rect 72292 1884 72298 1896
rect 72329 1887 72387 1893
rect 72329 1884 72341 1887
rect 72292 1856 72341 1884
rect 72292 1844 72298 1856
rect 72329 1853 72341 1856
rect 72375 1853 72387 1887
rect 72329 1847 72387 1853
rect 72973 1887 73031 1893
rect 72973 1853 72985 1887
rect 73019 1884 73031 1887
rect 73801 1887 73859 1893
rect 73801 1884 73813 1887
rect 73019 1856 73813 1884
rect 73019 1853 73031 1856
rect 72973 1847 73031 1853
rect 73801 1853 73813 1856
rect 73847 1853 73859 1887
rect 73801 1847 73859 1853
rect 55858 1816 55864 1828
rect 52840 1788 55864 1816
rect 55858 1776 55864 1788
rect 55916 1776 55922 1828
rect 60277 1819 60335 1825
rect 60277 1785 60289 1819
rect 60323 1816 60335 1819
rect 65794 1816 65800 1828
rect 60323 1788 65800 1816
rect 60323 1785 60335 1788
rect 60277 1779 60335 1785
rect 65794 1776 65800 1788
rect 65852 1776 65858 1828
rect 69382 1776 69388 1828
rect 69440 1776 69446 1828
rect 42567 1720 51948 1748
rect 56137 1751 56195 1757
rect 42567 1717 42579 1720
rect 42521 1711 42579 1717
rect 56137 1717 56149 1751
rect 56183 1748 56195 1751
rect 57238 1748 57244 1760
rect 56183 1720 57244 1748
rect 56183 1717 56195 1720
rect 56137 1711 56195 1717
rect 57238 1708 57244 1720
rect 57296 1708 57302 1760
rect 61105 1751 61163 1757
rect 61105 1717 61117 1751
rect 61151 1748 61163 1751
rect 62390 1748 62396 1760
rect 61151 1720 62396 1748
rect 61151 1717 61163 1720
rect 61105 1711 61163 1717
rect 62390 1708 62396 1720
rect 62448 1708 62454 1760
rect 64417 1751 64475 1757
rect 64417 1717 64429 1751
rect 64463 1748 64475 1751
rect 65150 1748 65156 1760
rect 64463 1720 65156 1748
rect 64463 1717 64475 1720
rect 64417 1711 64475 1717
rect 65150 1708 65156 1720
rect 65208 1708 65214 1760
rect 73154 1708 73160 1760
rect 73212 1748 73218 1760
rect 73249 1751 73307 1757
rect 73249 1748 73261 1751
rect 73212 1720 73261 1748
rect 73212 1708 73218 1720
rect 73249 1717 73261 1720
rect 73295 1717 73307 1751
rect 73249 1711 73307 1717
rect 1012 1658 74980 1680
rect 1012 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 74980 1658
rect 1012 1584 74980 1606
rect 22649 1547 22707 1553
rect 22649 1513 22661 1547
rect 22695 1544 22707 1547
rect 22922 1544 22928 1556
rect 22695 1516 22928 1544
rect 22695 1513 22707 1516
rect 22649 1507 22707 1513
rect 22922 1504 22928 1516
rect 22980 1504 22986 1556
rect 25225 1547 25283 1553
rect 25225 1513 25237 1547
rect 25271 1544 25283 1547
rect 26050 1544 26056 1556
rect 25271 1516 26056 1544
rect 25271 1513 25283 1516
rect 25225 1507 25283 1513
rect 26050 1504 26056 1516
rect 26108 1504 26114 1556
rect 27801 1547 27859 1553
rect 27801 1513 27813 1547
rect 27847 1544 27859 1547
rect 28626 1544 28632 1556
rect 27847 1516 28632 1544
rect 27847 1513 27859 1516
rect 27801 1507 27859 1513
rect 28626 1504 28632 1516
rect 28684 1504 28690 1556
rect 30377 1547 30435 1553
rect 30377 1513 30389 1547
rect 30423 1544 30435 1547
rect 31018 1544 31024 1556
rect 30423 1516 31024 1544
rect 30423 1513 30435 1516
rect 30377 1507 30435 1513
rect 31018 1504 31024 1516
rect 31076 1504 31082 1556
rect 32674 1504 32680 1556
rect 32732 1544 32738 1556
rect 37458 1544 37464 1556
rect 32732 1516 37464 1544
rect 32732 1504 32738 1516
rect 37458 1504 37464 1516
rect 37516 1504 37522 1556
rect 37550 1504 37556 1556
rect 37608 1544 37614 1556
rect 37921 1547 37979 1553
rect 37921 1544 37933 1547
rect 37608 1516 37933 1544
rect 37608 1504 37614 1516
rect 37921 1513 37933 1516
rect 37967 1513 37979 1547
rect 37921 1507 37979 1513
rect 41138 1504 41144 1556
rect 41196 1544 41202 1556
rect 41233 1547 41291 1553
rect 41233 1544 41245 1547
rect 41196 1516 41245 1544
rect 41196 1504 41202 1516
rect 41233 1513 41245 1516
rect 41279 1513 41291 1547
rect 41233 1507 41291 1513
rect 45370 1504 45376 1556
rect 45428 1504 45434 1556
rect 45554 1504 45560 1556
rect 45612 1544 45618 1556
rect 46385 1547 46443 1553
rect 46385 1544 46397 1547
rect 45612 1516 46397 1544
rect 45612 1504 45618 1516
rect 46385 1513 46397 1516
rect 46431 1513 46443 1547
rect 46385 1507 46443 1513
rect 47210 1504 47216 1556
rect 47268 1544 47274 1556
rect 48961 1547 49019 1553
rect 48961 1544 48973 1547
rect 47268 1516 48973 1544
rect 47268 1504 47274 1516
rect 48961 1513 48973 1516
rect 49007 1513 49019 1547
rect 48961 1507 49019 1513
rect 51258 1504 51264 1556
rect 51316 1544 51322 1556
rect 51537 1547 51595 1553
rect 51537 1544 51549 1547
rect 51316 1516 51549 1544
rect 51316 1504 51322 1516
rect 51537 1513 51549 1516
rect 51583 1513 51595 1547
rect 51537 1507 51595 1513
rect 61010 1504 61016 1556
rect 61068 1544 61074 1556
rect 61841 1547 61899 1553
rect 61841 1544 61853 1547
rect 61068 1516 61853 1544
rect 61068 1504 61074 1516
rect 61841 1513 61853 1516
rect 61887 1513 61899 1547
rect 61841 1507 61899 1513
rect 63862 1504 63868 1556
rect 63920 1544 63926 1556
rect 64417 1547 64475 1553
rect 64417 1544 64429 1547
rect 63920 1516 64429 1544
rect 63920 1504 63926 1516
rect 64417 1513 64429 1516
rect 64463 1513 64475 1547
rect 64417 1507 64475 1513
rect 69934 1504 69940 1556
rect 69992 1544 69998 1556
rect 70213 1547 70271 1553
rect 70213 1544 70225 1547
rect 69992 1516 70225 1544
rect 69992 1504 69998 1516
rect 70213 1513 70225 1516
rect 70259 1513 70271 1547
rect 70213 1507 70271 1513
rect 31110 1476 31116 1488
rect 22066 1448 31116 1476
rect 19150 1368 19156 1420
rect 19208 1408 19214 1420
rect 20254 1408 20260 1420
rect 19208 1380 20260 1408
rect 19208 1368 19214 1380
rect 20254 1368 20260 1380
rect 20312 1368 20318 1420
rect 20993 1411 21051 1417
rect 20993 1377 21005 1411
rect 21039 1408 21051 1411
rect 22066 1408 22094 1448
rect 31110 1436 31116 1448
rect 31168 1436 31174 1488
rect 31294 1436 31300 1488
rect 31352 1476 31358 1488
rect 41598 1476 41604 1488
rect 31352 1448 41604 1476
rect 31352 1436 31358 1448
rect 41598 1436 41604 1448
rect 41656 1436 41662 1488
rect 45388 1476 45416 1504
rect 47121 1479 47179 1485
rect 47121 1476 47133 1479
rect 45388 1448 47133 1476
rect 47121 1445 47133 1448
rect 47167 1445 47179 1479
rect 47121 1439 47179 1445
rect 21039 1380 22094 1408
rect 21039 1377 21051 1380
rect 20993 1371 21051 1377
rect 22830 1368 22836 1420
rect 22888 1408 22894 1420
rect 22888 1380 27200 1408
rect 22888 1368 22894 1380
rect 5074 1300 5080 1352
rect 5132 1300 5138 1352
rect 15286 1300 15292 1352
rect 15344 1340 15350 1352
rect 15381 1343 15439 1349
rect 15381 1340 15393 1343
rect 15344 1312 15393 1340
rect 15344 1300 15350 1312
rect 15381 1309 15393 1312
rect 15427 1309 15439 1343
rect 15381 1303 15439 1309
rect 15749 1343 15807 1349
rect 15749 1309 15761 1343
rect 15795 1340 15807 1343
rect 17494 1340 17500 1352
rect 15795 1312 17500 1340
rect 15795 1309 15807 1312
rect 15749 1303 15807 1309
rect 17494 1300 17500 1312
rect 17552 1300 17558 1352
rect 17770 1300 17776 1352
rect 17828 1300 17834 1352
rect 18049 1343 18107 1349
rect 18049 1340 18061 1343
rect 17880 1312 18061 1340
rect 3142 1232 3148 1284
rect 3200 1272 3206 1284
rect 3881 1275 3939 1281
rect 3881 1272 3893 1275
rect 3200 1244 3893 1272
rect 3200 1232 3206 1244
rect 3881 1241 3893 1244
rect 3927 1241 3939 1275
rect 3881 1235 3939 1241
rect 15838 1232 15844 1284
rect 15896 1272 15902 1284
rect 16761 1275 16819 1281
rect 16761 1272 16773 1275
rect 15896 1244 16773 1272
rect 15896 1232 15902 1244
rect 16761 1241 16773 1244
rect 16807 1241 16819 1275
rect 16761 1235 16819 1241
rect 15562 1164 15568 1216
rect 15620 1164 15626 1216
rect 16393 1207 16451 1213
rect 16393 1173 16405 1207
rect 16439 1204 16451 1207
rect 17880 1204 17908 1312
rect 18049 1309 18061 1312
rect 18095 1309 18107 1343
rect 18049 1303 18107 1309
rect 18325 1343 18383 1349
rect 18325 1309 18337 1343
rect 18371 1340 18383 1343
rect 19058 1340 19064 1352
rect 18371 1312 19064 1340
rect 18371 1309 18383 1312
rect 18325 1303 18383 1309
rect 19058 1300 19064 1312
rect 19116 1300 19122 1352
rect 19705 1343 19763 1349
rect 19705 1309 19717 1343
rect 19751 1309 19763 1343
rect 19705 1303 19763 1309
rect 19426 1232 19432 1284
rect 19484 1232 19490 1284
rect 19720 1272 19748 1303
rect 19794 1300 19800 1352
rect 19852 1300 19858 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22554 1340 22560 1352
rect 22051 1312 22560 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22554 1300 22560 1312
rect 22612 1300 22618 1352
rect 24121 1343 24179 1349
rect 24121 1309 24133 1343
rect 24167 1309 24179 1343
rect 24121 1303 24179 1309
rect 24673 1343 24731 1349
rect 24673 1309 24685 1343
rect 24719 1340 24731 1343
rect 26326 1340 26332 1352
rect 24719 1312 26332 1340
rect 24719 1309 24731 1312
rect 24673 1303 24731 1309
rect 22278 1272 22284 1284
rect 19720 1244 22284 1272
rect 22278 1232 22284 1244
rect 22336 1232 22342 1284
rect 23201 1275 23259 1281
rect 23201 1241 23213 1275
rect 23247 1272 23259 1275
rect 23566 1272 23572 1284
rect 23247 1244 23572 1272
rect 23247 1241 23259 1244
rect 23201 1235 23259 1241
rect 23566 1232 23572 1244
rect 23624 1232 23630 1284
rect 16439 1176 17908 1204
rect 24136 1204 24164 1303
rect 26326 1300 26332 1312
rect 26384 1300 26390 1352
rect 26697 1343 26755 1349
rect 26697 1309 26709 1343
rect 26743 1309 26755 1343
rect 26697 1303 26755 1309
rect 25774 1232 25780 1284
rect 25832 1232 25838 1284
rect 26510 1204 26516 1216
rect 24136 1176 26516 1204
rect 16439 1173 16451 1176
rect 16393 1167 16451 1173
rect 26510 1164 26516 1176
rect 26568 1164 26574 1216
rect 26712 1204 26740 1303
rect 27172 1272 27200 1380
rect 27982 1368 27988 1420
rect 28040 1408 28046 1420
rect 28353 1411 28411 1417
rect 28353 1408 28365 1411
rect 28040 1380 28365 1408
rect 28040 1368 28046 1380
rect 28353 1377 28365 1380
rect 28399 1377 28411 1411
rect 33042 1408 33048 1420
rect 28353 1371 28411 1377
rect 28460 1380 33048 1408
rect 27249 1343 27307 1349
rect 27249 1309 27261 1343
rect 27295 1340 27307 1343
rect 27798 1340 27804 1352
rect 27295 1312 27804 1340
rect 27295 1309 27307 1312
rect 27249 1303 27307 1309
rect 27798 1300 27804 1312
rect 27856 1300 27862 1352
rect 27893 1343 27951 1349
rect 27893 1309 27905 1343
rect 27939 1340 27951 1343
rect 27939 1336 28028 1340
rect 28074 1336 28080 1352
rect 27939 1312 28080 1336
rect 27939 1309 27951 1312
rect 27893 1303 27951 1309
rect 28000 1308 28080 1312
rect 28074 1300 28080 1308
rect 28132 1300 28138 1352
rect 28460 1272 28488 1380
rect 33042 1368 33048 1380
rect 33100 1368 33106 1420
rect 33152 1380 33364 1408
rect 28994 1300 29000 1352
rect 29052 1340 29058 1352
rect 29457 1343 29515 1349
rect 29457 1340 29469 1343
rect 29052 1312 29469 1340
rect 29052 1300 29058 1312
rect 29457 1309 29469 1312
rect 29503 1309 29515 1343
rect 29457 1303 29515 1309
rect 29825 1343 29883 1349
rect 29825 1309 29837 1343
rect 29871 1340 29883 1343
rect 30374 1340 30380 1352
rect 29871 1312 30380 1340
rect 29871 1309 29883 1312
rect 29825 1303 29883 1309
rect 30374 1300 30380 1312
rect 30432 1300 30438 1352
rect 30469 1343 30527 1349
rect 30469 1309 30481 1343
rect 30515 1309 30527 1343
rect 30469 1303 30527 1309
rect 32401 1343 32459 1349
rect 32401 1309 32413 1343
rect 32447 1340 32459 1343
rect 33152 1340 33180 1380
rect 32447 1312 33180 1340
rect 32447 1309 32459 1312
rect 32401 1303 32459 1309
rect 30484 1272 30512 1303
rect 33226 1300 33232 1352
rect 33284 1300 33290 1352
rect 33336 1340 33364 1380
rect 37918 1368 37924 1420
rect 37976 1408 37982 1420
rect 38473 1411 38531 1417
rect 38473 1408 38485 1411
rect 37976 1380 38485 1408
rect 37976 1368 37982 1380
rect 38473 1377 38485 1380
rect 38519 1377 38531 1411
rect 38473 1371 38531 1377
rect 41230 1368 41236 1420
rect 41288 1408 41294 1420
rect 42797 1411 42855 1417
rect 42797 1408 42809 1411
rect 41288 1380 42809 1408
rect 41288 1368 41294 1380
rect 42797 1377 42809 1380
rect 42843 1377 42855 1411
rect 42797 1371 42855 1377
rect 43070 1368 43076 1420
rect 43128 1408 43134 1420
rect 43128 1380 44404 1408
rect 43128 1368 43134 1380
rect 33502 1340 33508 1352
rect 33336 1312 33508 1340
rect 33502 1300 33508 1312
rect 33560 1300 33566 1352
rect 34977 1343 35035 1349
rect 34977 1309 34989 1343
rect 35023 1309 35035 1343
rect 34977 1303 35035 1309
rect 27172 1244 28488 1272
rect 29656 1244 30512 1272
rect 27890 1204 27896 1216
rect 26712 1176 27896 1204
rect 27890 1164 27896 1176
rect 27948 1164 27954 1216
rect 29656 1213 29684 1244
rect 31294 1232 31300 1284
rect 31352 1272 31358 1284
rect 31389 1275 31447 1281
rect 31389 1272 31401 1275
rect 31352 1244 31401 1272
rect 31352 1232 31358 1244
rect 31389 1241 31401 1244
rect 31435 1241 31447 1275
rect 31389 1235 31447 1241
rect 33134 1232 33140 1284
rect 33192 1272 33198 1284
rect 33965 1275 34023 1281
rect 33965 1272 33977 1275
rect 33192 1244 33977 1272
rect 33192 1232 33198 1244
rect 33965 1241 33977 1244
rect 34011 1241 34023 1275
rect 33965 1235 34023 1241
rect 29641 1207 29699 1213
rect 29641 1173 29653 1207
rect 29687 1173 29699 1207
rect 29641 1167 29699 1173
rect 32953 1207 33011 1213
rect 32953 1173 32965 1207
rect 32999 1204 33011 1207
rect 33594 1204 33600 1216
rect 32999 1176 33600 1204
rect 32999 1173 33011 1176
rect 32953 1167 33011 1173
rect 33594 1164 33600 1176
rect 33652 1164 33658 1216
rect 34992 1204 35020 1303
rect 35618 1300 35624 1352
rect 35676 1300 35682 1352
rect 37366 1300 37372 1352
rect 37424 1300 37430 1352
rect 37458 1300 37464 1352
rect 37516 1340 37522 1352
rect 38013 1343 38071 1349
rect 38013 1340 38025 1343
rect 37516 1312 38025 1340
rect 37516 1300 37522 1312
rect 38013 1309 38025 1312
rect 38059 1309 38071 1343
rect 38013 1303 38071 1309
rect 39758 1300 39764 1352
rect 39816 1300 39822 1352
rect 40770 1300 40776 1352
rect 40828 1340 40834 1352
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 40828 1312 41797 1340
rect 40828 1300 40834 1312
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41785 1303 41843 1309
rect 42426 1300 42432 1352
rect 42484 1300 42490 1352
rect 42886 1300 42892 1352
rect 42944 1340 42950 1352
rect 44376 1349 44404 1380
rect 44818 1368 44824 1420
rect 44876 1408 44882 1420
rect 45373 1411 45431 1417
rect 45373 1408 45385 1411
rect 44876 1380 45385 1408
rect 44876 1368 44882 1380
rect 45373 1377 45385 1380
rect 45419 1377 45431 1411
rect 45373 1371 45431 1377
rect 46198 1368 46204 1420
rect 46256 1408 46262 1420
rect 47949 1411 48007 1417
rect 47949 1408 47961 1411
rect 46256 1380 47961 1408
rect 46256 1368 46262 1380
rect 47949 1377 47961 1380
rect 47995 1377 48007 1411
rect 47949 1371 48007 1377
rect 49602 1368 49608 1420
rect 49660 1408 49666 1420
rect 50525 1411 50583 1417
rect 50525 1408 50537 1411
rect 49660 1380 50537 1408
rect 49660 1368 49666 1380
rect 50525 1377 50537 1380
rect 50571 1377 50583 1411
rect 50525 1371 50583 1377
rect 59446 1368 59452 1420
rect 59504 1408 59510 1420
rect 60829 1411 60887 1417
rect 60829 1408 60841 1411
rect 59504 1380 60841 1408
rect 59504 1368 59510 1380
rect 60829 1377 60841 1380
rect 60875 1377 60887 1411
rect 60829 1371 60887 1377
rect 62758 1368 62764 1420
rect 62816 1408 62822 1420
rect 63405 1411 63463 1417
rect 63405 1408 63417 1411
rect 62816 1380 63417 1408
rect 62816 1368 62822 1380
rect 63405 1377 63417 1380
rect 63451 1377 63463 1411
rect 63405 1371 63463 1377
rect 67726 1368 67732 1420
rect 67784 1408 67790 1420
rect 68557 1411 68615 1417
rect 68557 1408 68569 1411
rect 67784 1380 68569 1408
rect 67784 1368 67790 1380
rect 68557 1377 68569 1380
rect 68603 1377 68615 1411
rect 68557 1371 68615 1377
rect 71038 1368 71044 1420
rect 71096 1408 71102 1420
rect 71593 1411 71651 1417
rect 71593 1408 71605 1411
rect 71096 1380 71605 1408
rect 71096 1368 71102 1380
rect 71593 1377 71605 1380
rect 71639 1377 71651 1411
rect 71593 1371 71651 1377
rect 43809 1343 43867 1349
rect 43809 1340 43821 1343
rect 42944 1312 43821 1340
rect 42944 1300 42950 1312
rect 43809 1309 43821 1312
rect 43855 1309 43867 1343
rect 43809 1303 43867 1309
rect 44361 1343 44419 1349
rect 44361 1309 44373 1343
rect 44407 1309 44419 1343
rect 44361 1303 44419 1309
rect 44545 1343 44603 1349
rect 44545 1309 44557 1343
rect 44591 1340 44603 1343
rect 44726 1340 44732 1352
rect 44591 1312 44732 1340
rect 44591 1309 44603 1312
rect 44545 1303 44603 1309
rect 44726 1300 44732 1312
rect 44784 1300 44790 1352
rect 44910 1300 44916 1352
rect 44968 1300 44974 1352
rect 46937 1343 46995 1349
rect 46937 1340 46949 1343
rect 45020 1312 46949 1340
rect 35529 1275 35587 1281
rect 35529 1241 35541 1275
rect 35575 1272 35587 1275
rect 36170 1272 36176 1284
rect 35575 1244 36176 1272
rect 35575 1241 35587 1244
rect 35529 1235 35587 1241
rect 36170 1232 36176 1244
rect 36228 1232 36234 1284
rect 36262 1232 36268 1284
rect 36320 1272 36326 1284
rect 36541 1275 36599 1281
rect 36541 1272 36553 1275
rect 36320 1244 36553 1272
rect 36320 1232 36326 1244
rect 36541 1241 36553 1244
rect 36587 1241 36599 1275
rect 36541 1235 36599 1241
rect 39574 1232 39580 1284
rect 39632 1272 39638 1284
rect 40681 1275 40739 1281
rect 40681 1272 40693 1275
rect 39632 1244 40693 1272
rect 39632 1232 39638 1244
rect 40681 1241 40693 1244
rect 40727 1241 40739 1275
rect 40681 1235 40739 1241
rect 43990 1232 43996 1284
rect 44048 1272 44054 1284
rect 45020 1272 45048 1312
rect 46937 1309 46949 1312
rect 46983 1309 46995 1343
rect 46937 1303 46995 1309
rect 47305 1343 47363 1349
rect 47305 1309 47317 1343
rect 47351 1309 47363 1343
rect 47305 1303 47363 1309
rect 44048 1244 45048 1272
rect 44048 1232 44054 1244
rect 45094 1232 45100 1284
rect 45152 1272 45158 1284
rect 47320 1272 47348 1303
rect 47394 1300 47400 1352
rect 47452 1340 47458 1352
rect 47489 1343 47547 1349
rect 47489 1340 47501 1343
rect 47452 1312 47501 1340
rect 47452 1300 47458 1312
rect 47489 1309 47501 1312
rect 47535 1309 47547 1343
rect 47489 1303 47547 1309
rect 49418 1300 49424 1352
rect 49476 1340 49482 1352
rect 49513 1343 49571 1349
rect 49513 1340 49525 1343
rect 49476 1312 49525 1340
rect 49476 1300 49482 1312
rect 49513 1309 49525 1312
rect 49559 1309 49571 1343
rect 49513 1303 49571 1309
rect 50062 1300 50068 1352
rect 50120 1300 50126 1352
rect 50614 1300 50620 1352
rect 50672 1340 50678 1352
rect 52089 1343 52147 1349
rect 52089 1340 52101 1343
rect 50672 1312 52101 1340
rect 50672 1300 50678 1312
rect 52089 1309 52101 1312
rect 52135 1309 52147 1343
rect 52089 1303 52147 1309
rect 52638 1300 52644 1352
rect 52696 1300 52702 1352
rect 53834 1300 53840 1352
rect 53892 1340 53898 1352
rect 54113 1343 54171 1349
rect 54113 1340 54125 1343
rect 53892 1312 54125 1340
rect 53892 1300 53898 1312
rect 54113 1309 54125 1312
rect 54159 1309 54171 1343
rect 54665 1343 54723 1349
rect 54665 1340 54677 1343
rect 54113 1303 54171 1309
rect 54220 1312 54677 1340
rect 45152 1244 47348 1272
rect 45152 1232 45158 1244
rect 51166 1232 51172 1284
rect 51224 1272 51230 1284
rect 53561 1275 53619 1281
rect 53561 1272 53573 1275
rect 51224 1244 53573 1272
rect 51224 1232 51230 1244
rect 53561 1241 53573 1244
rect 53607 1241 53619 1275
rect 53561 1235 53619 1241
rect 35710 1204 35716 1216
rect 34992 1176 35716 1204
rect 35710 1164 35716 1176
rect 35768 1164 35774 1216
rect 44729 1207 44787 1213
rect 44729 1173 44741 1207
rect 44775 1204 44787 1207
rect 46014 1204 46020 1216
rect 44775 1176 46020 1204
rect 44775 1173 44787 1176
rect 44729 1167 44787 1173
rect 46014 1164 46020 1176
rect 46072 1164 46078 1216
rect 52270 1164 52276 1216
rect 52328 1204 52334 1216
rect 54220 1204 54248 1312
rect 54665 1309 54677 1312
rect 54711 1309 54723 1343
rect 54665 1303 54723 1309
rect 55214 1300 55220 1352
rect 55272 1300 55278 1352
rect 56686 1300 56692 1352
rect 56744 1300 56750 1352
rect 57238 1300 57244 1352
rect 57296 1300 57302 1352
rect 57974 1300 57980 1352
rect 58032 1300 58038 1352
rect 59354 1300 59360 1352
rect 59412 1300 59418 1352
rect 59909 1343 59967 1349
rect 59909 1309 59921 1343
rect 59955 1309 59967 1343
rect 59909 1303 59967 1309
rect 54570 1232 54576 1284
rect 54628 1272 54634 1284
rect 56137 1275 56195 1281
rect 56137 1272 56149 1275
rect 54628 1244 56149 1272
rect 54628 1232 54634 1244
rect 56137 1241 56149 1244
rect 56183 1241 56195 1275
rect 56137 1235 56195 1241
rect 57790 1232 57796 1284
rect 57848 1272 57854 1284
rect 58805 1275 58863 1281
rect 58805 1272 58817 1275
rect 57848 1244 58817 1272
rect 57848 1232 57854 1244
rect 58805 1241 58817 1244
rect 58851 1241 58863 1275
rect 58805 1235 58863 1241
rect 58894 1232 58900 1284
rect 58952 1272 58958 1284
rect 59924 1272 59952 1303
rect 60366 1300 60372 1352
rect 60424 1300 60430 1352
rect 62390 1300 62396 1352
rect 62448 1300 62454 1352
rect 63034 1300 63040 1352
rect 63092 1300 63098 1352
rect 63862 1300 63868 1352
rect 63920 1340 63926 1352
rect 64969 1343 65027 1349
rect 64969 1340 64981 1343
rect 63920 1312 64981 1340
rect 63920 1300 63926 1312
rect 64969 1309 64981 1312
rect 65015 1309 65027 1343
rect 64969 1303 65027 1309
rect 65150 1300 65156 1352
rect 65208 1340 65214 1352
rect 65521 1343 65579 1349
rect 65521 1340 65533 1343
rect 65208 1312 65533 1340
rect 65208 1300 65214 1312
rect 65521 1309 65533 1312
rect 65567 1309 65579 1343
rect 65521 1303 65579 1309
rect 66254 1300 66260 1352
rect 66312 1300 66318 1352
rect 68278 1300 68284 1352
rect 68336 1300 68342 1352
rect 68830 1300 68836 1352
rect 68888 1340 68894 1352
rect 69569 1343 69627 1349
rect 69569 1340 69581 1343
rect 68888 1312 69581 1340
rect 68888 1300 68894 1312
rect 69569 1309 69581 1312
rect 69615 1309 69627 1343
rect 69569 1303 69627 1309
rect 71222 1300 71228 1352
rect 71280 1300 71286 1352
rect 73065 1343 73123 1349
rect 73065 1309 73077 1343
rect 73111 1340 73123 1343
rect 73154 1340 73160 1352
rect 73111 1312 73160 1340
rect 73111 1309 73123 1312
rect 73065 1303 73123 1309
rect 73154 1300 73160 1312
rect 73212 1300 73218 1352
rect 73246 1300 73252 1352
rect 73304 1300 73310 1352
rect 58952 1244 59952 1272
rect 65797 1275 65855 1281
rect 58952 1232 58958 1244
rect 65797 1241 65809 1275
rect 65843 1241 65855 1275
rect 65797 1235 65855 1241
rect 52328 1176 54248 1204
rect 65812 1204 65840 1235
rect 66070 1232 66076 1284
rect 66128 1272 66134 1284
rect 67085 1275 67143 1281
rect 67085 1272 67097 1275
rect 66128 1244 67097 1272
rect 66128 1232 66134 1244
rect 67085 1241 67097 1244
rect 67131 1241 67143 1275
rect 67085 1235 67143 1241
rect 70026 1232 70032 1284
rect 70084 1272 70090 1284
rect 72789 1275 72847 1281
rect 72789 1272 72801 1275
rect 70084 1244 72801 1272
rect 70084 1232 70090 1244
rect 72789 1241 72801 1244
rect 72835 1241 72847 1275
rect 72789 1235 72847 1241
rect 74169 1275 74227 1281
rect 74169 1241 74181 1275
rect 74215 1241 74227 1275
rect 74169 1235 74227 1241
rect 67358 1204 67364 1216
rect 65812 1176 67364 1204
rect 52328 1164 52334 1176
rect 67358 1164 67364 1176
rect 67416 1164 67422 1216
rect 72694 1164 72700 1216
rect 72752 1204 72758 1216
rect 74184 1204 74212 1235
rect 72752 1176 74212 1204
rect 72752 1164 72758 1176
rect 1012 1114 74980 1136
rect 1012 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74980 1114
rect 1012 1040 74980 1062
rect 5074 960 5080 1012
rect 5132 1000 5138 1012
rect 23934 1000 23940 1012
rect 5132 972 23940 1000
rect 5132 960 5138 972
rect 23934 960 23940 972
rect 23992 960 23998 1012
rect 31386 960 31392 1012
rect 31444 1000 31450 1012
rect 35618 1000 35624 1012
rect 31444 972 35624 1000
rect 31444 960 31450 972
rect 35618 960 35624 972
rect 35676 960 35682 1012
rect 15562 892 15568 944
rect 15620 932 15626 944
rect 20714 932 20720 944
rect 15620 904 20720 932
rect 15620 892 15626 904
rect 20714 892 20720 904
rect 20772 892 20778 944
rect 27798 892 27804 944
rect 27856 932 27862 944
rect 28534 932 28540 944
rect 27856 904 28540 932
rect 27856 892 27862 904
rect 28534 892 28540 904
rect 28592 892 28598 944
rect 19426 824 19432 876
rect 19484 864 19490 876
rect 43622 864 43628 876
rect 19484 836 43628 864
rect 19484 824 19490 836
rect 43622 824 43628 836
rect 43680 824 43686 876
<< via1 >>
rect 74210 85926 74262 85978
rect 74274 85926 74326 85978
rect 74338 85926 74390 85978
rect 74402 85926 74454 85978
rect 74466 85926 74518 85978
rect 71858 85382 71910 85434
rect 71922 85382 71974 85434
rect 71986 85382 72038 85434
rect 72050 85382 72102 85434
rect 72114 85382 72166 85434
rect 74210 84838 74262 84890
rect 74274 84838 74326 84890
rect 74338 84838 74390 84890
rect 74402 84838 74454 84890
rect 74466 84838 74518 84890
rect 71858 84294 71910 84346
rect 71922 84294 71974 84346
rect 71986 84294 72038 84346
rect 72050 84294 72102 84346
rect 72114 84294 72166 84346
rect 64880 84192 64932 84244
rect 74210 83750 74262 83802
rect 74274 83750 74326 83802
rect 74338 83750 74390 83802
rect 74402 83750 74454 83802
rect 74466 83750 74518 83802
rect 71858 83206 71910 83258
rect 71922 83206 71974 83258
rect 71986 83206 72038 83258
rect 72050 83206 72102 83258
rect 72114 83206 72166 83258
rect 66996 83104 67048 83156
rect 69664 82968 69716 83020
rect 74210 82662 74262 82714
rect 74274 82662 74326 82714
rect 74338 82662 74390 82714
rect 74402 82662 74454 82714
rect 74466 82662 74518 82714
rect 71858 82118 71910 82170
rect 71922 82118 71974 82170
rect 71986 82118 72038 82170
rect 72050 82118 72102 82170
rect 72114 82118 72166 82170
rect 64880 81744 64932 81796
rect 74210 81574 74262 81626
rect 74274 81574 74326 81626
rect 74338 81574 74390 81626
rect 74402 81574 74454 81626
rect 74466 81574 74518 81626
rect 71858 81030 71910 81082
rect 71922 81030 71974 81082
rect 71986 81030 72038 81082
rect 72050 81030 72102 81082
rect 72114 81030 72166 81082
rect 67088 80928 67140 80980
rect 69756 80792 69808 80844
rect 74210 80486 74262 80538
rect 74274 80486 74326 80538
rect 74338 80486 74390 80538
rect 74402 80486 74454 80538
rect 74466 80486 74518 80538
rect 71858 79942 71910 79994
rect 71922 79942 71974 79994
rect 71986 79942 72038 79994
rect 72050 79942 72102 79994
rect 72114 79942 72166 79994
rect 64880 79840 64932 79892
rect 74210 79398 74262 79450
rect 74274 79398 74326 79450
rect 74338 79398 74390 79450
rect 74402 79398 74454 79450
rect 74466 79398 74518 79450
rect 71858 78854 71910 78906
rect 71922 78854 71974 78906
rect 71986 78854 72038 78906
rect 72050 78854 72102 78906
rect 72114 78854 72166 78906
rect 66444 78684 66496 78736
rect 69940 78616 69992 78668
rect 74210 78310 74262 78362
rect 74274 78310 74326 78362
rect 74338 78310 74390 78362
rect 74402 78310 74454 78362
rect 74466 78310 74518 78362
rect 71858 77766 71910 77818
rect 71922 77766 71974 77818
rect 71986 77766 72038 77818
rect 72050 77766 72102 77818
rect 72114 77766 72166 77818
rect 64880 77664 64932 77716
rect 74210 77222 74262 77274
rect 74274 77222 74326 77274
rect 74338 77222 74390 77274
rect 74402 77222 74454 77274
rect 74466 77222 74518 77274
rect 71858 76678 71910 76730
rect 71922 76678 71974 76730
rect 71986 76678 72038 76730
rect 72050 76678 72102 76730
rect 72114 76678 72166 76730
rect 66260 76508 66312 76560
rect 68468 76440 68520 76492
rect 74210 76134 74262 76186
rect 74274 76134 74326 76186
rect 74338 76134 74390 76186
rect 74402 76134 74454 76186
rect 74466 76134 74518 76186
rect 71858 75590 71910 75642
rect 71922 75590 71974 75642
rect 71986 75590 72038 75642
rect 72050 75590 72102 75642
rect 72114 75590 72166 75642
rect 64880 75148 64932 75200
rect 74210 75046 74262 75098
rect 74274 75046 74326 75098
rect 74338 75046 74390 75098
rect 74402 75046 74454 75098
rect 74466 75046 74518 75098
rect 67640 74604 67692 74656
rect 71858 74502 71910 74554
rect 71922 74502 71974 74554
rect 71986 74502 72038 74554
rect 72050 74502 72102 74554
rect 72114 74502 72166 74554
rect 66168 74060 66220 74112
rect 74210 73958 74262 74010
rect 74274 73958 74326 74010
rect 74338 73958 74390 74010
rect 74402 73958 74454 74010
rect 74466 73958 74518 74010
rect 71858 73414 71910 73466
rect 71922 73414 71974 73466
rect 71986 73414 72038 73466
rect 72050 73414 72102 73466
rect 72114 73414 72166 73466
rect 64880 73176 64932 73228
rect 74210 72870 74262 72922
rect 74274 72870 74326 72922
rect 74338 72870 74390 72922
rect 74402 72870 74454 72922
rect 74466 72870 74518 72922
rect 71858 72326 71910 72378
rect 71922 72326 71974 72378
rect 71986 72326 72038 72378
rect 72050 72326 72102 72378
rect 72114 72326 72166 72378
rect 66352 72156 66404 72208
rect 65984 71884 66036 71936
rect 74210 71782 74262 71834
rect 74274 71782 74326 71834
rect 74338 71782 74390 71834
rect 74402 71782 74454 71834
rect 74466 71782 74518 71834
rect 71858 71238 71910 71290
rect 71922 71238 71974 71290
rect 71986 71238 72038 71290
rect 72050 71238 72102 71290
rect 72114 71238 72166 71290
rect 64880 71068 64932 71120
rect 74210 70694 74262 70746
rect 74274 70694 74326 70746
rect 74338 70694 74390 70746
rect 74402 70694 74454 70746
rect 74466 70694 74518 70746
rect 71858 70150 71910 70202
rect 71922 70150 71974 70202
rect 71986 70150 72038 70202
rect 72050 70150 72102 70202
rect 72114 70150 72166 70202
rect 65524 69980 65576 70032
rect 63684 69572 63736 69624
rect 74210 69606 74262 69658
rect 74274 69606 74326 69658
rect 74338 69606 74390 69658
rect 74402 69606 74454 69658
rect 74466 69606 74518 69658
rect 71858 69062 71910 69114
rect 71922 69062 71974 69114
rect 71986 69062 72038 69114
rect 72050 69062 72102 69114
rect 72114 69062 72166 69114
rect 64880 68960 64932 69012
rect 66536 68960 66588 69012
rect 74210 68518 74262 68570
rect 74274 68518 74326 68570
rect 74338 68518 74390 68570
rect 74402 68518 74454 68570
rect 74466 68518 74518 68570
rect 71858 67974 71910 68026
rect 71922 67974 71974 68026
rect 71986 67974 72038 68026
rect 72050 67974 72102 68026
rect 72114 67974 72166 68026
rect 65892 67804 65944 67856
rect 64604 67600 64656 67652
rect 74210 67430 74262 67482
rect 74274 67430 74326 67482
rect 74338 67430 74390 67482
rect 74402 67430 74454 67482
rect 74466 67430 74518 67482
rect 71858 66886 71910 66938
rect 71922 66886 71974 66938
rect 71986 66886 72038 66938
rect 72050 66886 72102 66938
rect 72114 66886 72166 66938
rect 64880 66444 64932 66496
rect 74210 66342 74262 66394
rect 74274 66342 74326 66394
rect 74338 66342 74390 66394
rect 74402 66342 74454 66394
rect 74466 66342 74518 66394
rect 71858 65798 71910 65850
rect 71922 65798 71974 65850
rect 71986 65798 72038 65850
rect 72050 65798 72102 65850
rect 72114 65798 72166 65850
rect 65432 65628 65484 65680
rect 65708 65356 65760 65408
rect 74210 65254 74262 65306
rect 74274 65254 74326 65306
rect 74338 65254 74390 65306
rect 74402 65254 74454 65306
rect 74466 65254 74518 65306
rect 71858 64710 71910 64762
rect 71922 64710 71974 64762
rect 71986 64710 72038 64762
rect 72050 64710 72102 64762
rect 72114 64710 72166 64762
rect 64880 64268 64932 64320
rect 74210 64166 74262 64218
rect 74274 64166 74326 64218
rect 74338 64166 74390 64218
rect 74402 64166 74454 64218
rect 74466 64166 74518 64218
rect 71858 63622 71910 63674
rect 71922 63622 71974 63674
rect 71986 63622 72038 63674
rect 72050 63622 72102 63674
rect 72114 63622 72166 63674
rect 65340 63520 65392 63572
rect 69020 63384 69072 63436
rect 74210 63078 74262 63130
rect 74274 63078 74326 63130
rect 74338 63078 74390 63130
rect 74402 63078 74454 63130
rect 74466 63078 74518 63130
rect 71858 62534 71910 62586
rect 71922 62534 71974 62586
rect 71986 62534 72038 62586
rect 72050 62534 72102 62586
rect 72114 62534 72166 62586
rect 64880 62092 64932 62144
rect 74210 61990 74262 62042
rect 74274 61990 74326 62042
rect 74338 61990 74390 62042
rect 74402 61990 74454 62042
rect 74466 61990 74518 62042
rect 71858 61446 71910 61498
rect 71922 61446 71974 61498
rect 71986 61446 72038 61498
rect 72050 61446 72102 61498
rect 72114 61446 72166 61498
rect 65248 61276 65300 61328
rect 63592 60868 63644 60920
rect 74210 60902 74262 60954
rect 74274 60902 74326 60954
rect 74338 60902 74390 60954
rect 74402 60902 74454 60954
rect 74466 60902 74518 60954
rect 71858 60358 71910 60410
rect 71922 60358 71974 60410
rect 71986 60358 72038 60410
rect 72050 60358 72102 60410
rect 72114 60358 72166 60410
rect 64880 60188 64932 60240
rect 74210 59814 74262 59866
rect 74274 59814 74326 59866
rect 74338 59814 74390 59866
rect 74402 59814 74454 59866
rect 74466 59814 74518 59866
rect 71858 59270 71910 59322
rect 71922 59270 71974 59322
rect 71986 59270 72038 59322
rect 72050 59270 72102 59322
rect 72114 59270 72166 59322
rect 65156 59100 65208 59152
rect 70768 59032 70820 59084
rect 74210 58726 74262 58778
rect 74274 58726 74326 58778
rect 74338 58726 74390 58778
rect 74402 58726 74454 58778
rect 74466 58726 74518 58778
rect 71858 58182 71910 58234
rect 71922 58182 71974 58234
rect 71986 58182 72038 58234
rect 72050 58182 72102 58234
rect 72114 58182 72166 58234
rect 64880 58012 64932 58064
rect 74210 57638 74262 57690
rect 74274 57638 74326 57690
rect 74338 57638 74390 57690
rect 74402 57638 74454 57690
rect 74466 57638 74518 57690
rect 71858 57094 71910 57146
rect 71922 57094 71974 57146
rect 71986 57094 72038 57146
rect 72050 57094 72102 57146
rect 72114 57094 72166 57146
rect 68100 56992 68152 57044
rect 65800 56652 65852 56704
rect 74210 56550 74262 56602
rect 74274 56550 74326 56602
rect 74338 56550 74390 56602
rect 74402 56550 74454 56602
rect 74466 56550 74518 56602
rect 71858 56006 71910 56058
rect 71922 56006 71974 56058
rect 71986 56006 72038 56058
rect 72050 56006 72102 56058
rect 72114 56006 72166 56058
rect 64880 55564 64932 55616
rect 74210 55462 74262 55514
rect 74274 55462 74326 55514
rect 74338 55462 74390 55514
rect 74402 55462 74454 55514
rect 74466 55462 74518 55514
rect 71858 54918 71910 54970
rect 71922 54918 71974 54970
rect 71986 54918 72038 54970
rect 72050 54918 72102 54970
rect 72114 54918 72166 54970
rect 67548 54748 67600 54800
rect 69112 54612 69164 54664
rect 74210 54374 74262 54426
rect 74274 54374 74326 54426
rect 74338 54374 74390 54426
rect 74402 54374 74454 54426
rect 74466 54374 74518 54426
rect 71858 53830 71910 53882
rect 71922 53830 71974 53882
rect 71986 53830 72038 53882
rect 72050 53830 72102 53882
rect 72114 53830 72166 53882
rect 64880 53524 64932 53576
rect 74210 53286 74262 53338
rect 74274 53286 74326 53338
rect 74338 53286 74390 53338
rect 74402 53286 74454 53338
rect 74466 53286 74518 53338
rect 66904 53116 66956 53168
rect 71858 52742 71910 52794
rect 71922 52742 71974 52794
rect 71986 52742 72038 52794
rect 72050 52742 72102 52794
rect 72114 52742 72166 52794
rect 68192 52640 68244 52692
rect 63500 52572 63552 52624
rect 65616 52479 65668 52488
rect 65616 52445 65625 52479
rect 65625 52445 65659 52479
rect 65659 52445 65668 52479
rect 65616 52436 65668 52445
rect 74210 52198 74262 52250
rect 74274 52198 74326 52250
rect 74338 52198 74390 52250
rect 74402 52198 74454 52250
rect 74466 52198 74518 52250
rect 65616 52096 65668 52148
rect 71858 51654 71910 51706
rect 71922 51654 71974 51706
rect 71986 51654 72038 51706
rect 72050 51654 72102 51706
rect 72114 51654 72166 51706
rect 64880 51484 64932 51536
rect 66628 51484 66680 51536
rect 74210 51110 74262 51162
rect 74274 51110 74326 51162
rect 74338 51110 74390 51162
rect 74402 51110 74454 51162
rect 74466 51110 74518 51162
rect 71858 50566 71910 50618
rect 71922 50566 71974 50618
rect 71986 50566 72038 50618
rect 72050 50566 72102 50618
rect 72114 50566 72166 50618
rect 67364 50396 67416 50448
rect 63500 50260 63552 50312
rect 74210 50022 74262 50074
rect 74274 50022 74326 50074
rect 74338 50022 74390 50074
rect 74402 50022 74454 50074
rect 74466 50022 74518 50074
rect 71858 49478 71910 49530
rect 71922 49478 71974 49530
rect 71986 49478 72038 49530
rect 72050 49478 72102 49530
rect 72114 49478 72166 49530
rect 63408 48769 63460 48821
rect 74210 48934 74262 48986
rect 74274 48934 74326 48986
rect 74338 48934 74390 48986
rect 74402 48934 74454 48986
rect 74466 48934 74518 48986
rect 71858 48390 71910 48442
rect 71922 48390 71974 48442
rect 71986 48390 72038 48442
rect 72050 48390 72102 48442
rect 72114 48390 72166 48442
rect 63500 48061 63552 48113
rect 74210 47846 74262 47898
rect 74274 47846 74326 47898
rect 74338 47846 74390 47898
rect 74402 47846 74454 47898
rect 74466 47846 74518 47898
rect 63868 47676 63920 47728
rect 68560 47472 68612 47524
rect 71858 47302 71910 47354
rect 71922 47302 71974 47354
rect 71986 47302 72038 47354
rect 72050 47302 72102 47354
rect 72114 47302 72166 47354
rect 64788 46996 64840 47048
rect 67180 46996 67232 47048
rect 66812 46928 66864 46980
rect 74210 46758 74262 46810
rect 74274 46758 74326 46810
rect 74338 46758 74390 46810
rect 74402 46758 74454 46810
rect 74466 46758 74518 46810
rect 71858 46214 71910 46266
rect 71922 46214 71974 46266
rect 71986 46214 72038 46266
rect 72050 46214 72102 46266
rect 72114 46214 72166 46266
rect 68376 45976 68428 46028
rect 63960 45704 64012 45756
rect 74210 45670 74262 45722
rect 74274 45670 74326 45722
rect 74338 45670 74390 45722
rect 74402 45670 74454 45722
rect 74466 45670 74518 45722
rect 63868 45228 63920 45280
rect 71858 45126 71910 45178
rect 71922 45126 71974 45178
rect 71986 45126 72038 45178
rect 72050 45126 72102 45178
rect 72114 45126 72166 45178
rect 64880 44820 64932 44872
rect 74210 44582 74262 44634
rect 74274 44582 74326 44634
rect 74338 44582 74390 44634
rect 74402 44582 74454 44634
rect 74466 44582 74518 44634
rect 68284 44480 68336 44532
rect 67732 44412 67784 44464
rect 71858 44038 71910 44090
rect 71922 44038 71974 44090
rect 71986 44038 72038 44090
rect 72050 44038 72102 44090
rect 72114 44038 72166 44090
rect 64052 43800 64104 43852
rect 74210 43494 74262 43546
rect 74274 43494 74326 43546
rect 74338 43494 74390 43546
rect 74402 43494 74454 43546
rect 74466 43494 74518 43546
rect 70492 43256 70544 43308
rect 68744 43052 68796 43104
rect 71858 42950 71910 43002
rect 71922 42950 71974 43002
rect 71986 42950 72038 43002
rect 72050 42950 72102 43002
rect 72114 42950 72166 43002
rect 66996 42712 67048 42764
rect 70032 42644 70084 42696
rect 74210 42406 74262 42458
rect 74274 42406 74326 42458
rect 74338 42406 74390 42458
rect 74402 42406 74454 42458
rect 74466 42406 74518 42458
rect 71858 41862 71910 41914
rect 71922 41862 71974 41914
rect 71986 41862 72038 41914
rect 72050 41862 72102 41914
rect 72114 41862 72166 41914
rect 67088 41803 67140 41812
rect 67088 41769 67097 41803
rect 67097 41769 67131 41803
rect 67131 41769 67140 41803
rect 67088 41760 67140 41769
rect 65064 41692 65116 41744
rect 70124 41556 70176 41608
rect 74210 41318 74262 41370
rect 74274 41318 74326 41370
rect 74338 41318 74390 41370
rect 74402 41318 74454 41370
rect 74466 41318 74518 41370
rect 64972 40944 65024 40996
rect 67916 40876 67968 40928
rect 71858 40774 71910 40826
rect 71922 40774 71974 40826
rect 71986 40774 72038 40826
rect 72050 40774 72102 40826
rect 72114 40774 72166 40826
rect 66444 40715 66496 40724
rect 66444 40681 66453 40715
rect 66453 40681 66487 40715
rect 66487 40681 66496 40715
rect 66444 40672 66496 40681
rect 69204 40468 69256 40520
rect 74210 40230 74262 40282
rect 74274 40230 74326 40282
rect 74338 40230 74390 40282
rect 74402 40230 74454 40282
rect 74466 40230 74518 40282
rect 65064 39788 65116 39840
rect 71858 39686 71910 39738
rect 71922 39686 71974 39738
rect 71986 39686 72038 39738
rect 72050 39686 72102 39738
rect 72114 39686 72166 39738
rect 66260 39584 66312 39636
rect 67456 39380 67508 39432
rect 74210 39142 74262 39194
rect 74274 39142 74326 39194
rect 74338 39142 74390 39194
rect 74402 39142 74454 39194
rect 74466 39142 74518 39194
rect 64972 38836 65024 38888
rect 68008 38700 68060 38752
rect 71858 38598 71910 38650
rect 71922 38598 71974 38650
rect 71986 38598 72038 38650
rect 72050 38598 72102 38650
rect 72114 38598 72166 38650
rect 67640 38496 67692 38548
rect 66996 38292 67048 38344
rect 74210 38054 74262 38106
rect 74274 38054 74326 38106
rect 74338 38054 74390 38106
rect 74402 38054 74454 38106
rect 74466 38054 74518 38106
rect 71858 37510 71910 37562
rect 71922 37510 71974 37562
rect 71986 37510 72038 37562
rect 72050 37510 72102 37562
rect 72114 37510 72166 37562
rect 65064 37340 65116 37392
rect 67272 37204 67324 37256
rect 66352 37136 66404 37188
rect 74210 36966 74262 37018
rect 74274 36966 74326 37018
rect 74338 36966 74390 37018
rect 74402 36966 74454 37018
rect 74466 36966 74518 37018
rect 66076 36524 66128 36576
rect 71858 36422 71910 36474
rect 71922 36422 71974 36474
rect 71986 36422 72038 36474
rect 72050 36422 72102 36474
rect 72114 36422 72166 36474
rect 65524 36320 65576 36372
rect 69296 36252 69348 36304
rect 66352 36116 66404 36168
rect 74210 35878 74262 35930
rect 74274 35878 74326 35930
rect 74338 35878 74390 35930
rect 74402 35878 74454 35930
rect 74466 35878 74518 35930
rect 66536 35751 66588 35760
rect 66536 35717 66545 35751
rect 66545 35717 66579 35751
rect 66579 35717 66588 35751
rect 66536 35708 66588 35717
rect 70584 35640 70636 35692
rect 71858 35334 71910 35386
rect 71922 35334 71974 35386
rect 71986 35334 72038 35386
rect 72050 35334 72102 35386
rect 72114 35334 72166 35386
rect 65892 35232 65944 35284
rect 64880 35164 64932 35216
rect 65064 35164 65116 35216
rect 67088 35028 67140 35080
rect 74210 34790 74262 34842
rect 74274 34790 74326 34842
rect 74338 34790 74390 34842
rect 74402 34790 74454 34842
rect 74466 34790 74518 34842
rect 65524 34552 65576 34604
rect 71858 34246 71910 34298
rect 71922 34246 71974 34298
rect 71986 34246 72038 34298
rect 72050 34246 72102 34298
rect 72114 34246 72166 34298
rect 66904 34187 66956 34196
rect 66904 34153 66913 34187
rect 66913 34153 66947 34187
rect 66947 34153 66956 34187
rect 66904 34144 66956 34153
rect 64696 33940 64748 33992
rect 65616 33915 65668 33924
rect 65616 33881 65625 33915
rect 65625 33881 65659 33915
rect 65659 33881 65668 33915
rect 65616 33872 65668 33881
rect 74210 33702 74262 33754
rect 74274 33702 74326 33754
rect 74338 33702 74390 33754
rect 74402 33702 74454 33754
rect 74466 33702 74518 33754
rect 65432 33600 65484 33652
rect 66720 33396 66772 33448
rect 64880 33260 64932 33312
rect 71858 33158 71910 33210
rect 71922 33158 71974 33210
rect 71986 33158 72038 33210
rect 72050 33158 72102 33210
rect 72114 33158 72166 33210
rect 65340 33056 65392 33108
rect 66444 32852 66496 32904
rect 74210 32614 74262 32666
rect 74274 32614 74326 32666
rect 74338 32614 74390 32666
rect 74402 32614 74454 32666
rect 74466 32614 74518 32666
rect 65248 32172 65300 32224
rect 63500 32092 63552 32144
rect 71858 32070 71910 32122
rect 71922 32070 71974 32122
rect 71986 32070 72038 32122
rect 72050 32070 72102 32122
rect 72114 32070 72166 32122
rect 65340 31968 65392 32020
rect 66260 31807 66312 31816
rect 66260 31773 66269 31807
rect 66269 31773 66303 31807
rect 66303 31773 66312 31807
rect 66260 31764 66312 31773
rect 74210 31526 74262 31578
rect 74274 31526 74326 31578
rect 74338 31526 74390 31578
rect 74402 31526 74454 31578
rect 74466 31526 74518 31578
rect 64880 31084 64932 31136
rect 71858 30982 71910 31034
rect 71922 30982 71974 31034
rect 71986 30982 72038 31034
rect 72050 30982 72102 31034
rect 72114 30982 72166 31034
rect 65156 30880 65208 30932
rect 66536 30676 66588 30728
rect 74210 30438 74262 30490
rect 74274 30438 74326 30490
rect 74338 30438 74390 30490
rect 74402 30438 74454 30490
rect 74466 30438 74518 30490
rect 65340 29996 65392 30048
rect 71858 29894 71910 29946
rect 71922 29894 71974 29946
rect 71986 29894 72038 29946
rect 72050 29894 72102 29946
rect 72114 29894 72166 29946
rect 68100 29792 68152 29844
rect 63776 29588 63828 29640
rect 66996 29588 67048 29640
rect 74210 29350 74262 29402
rect 74274 29350 74326 29402
rect 74338 29350 74390 29402
rect 74402 29350 74454 29402
rect 74466 29350 74518 29402
rect 71858 28806 71910 28858
rect 71922 28806 71974 28858
rect 71986 28806 72038 28858
rect 72050 28806 72102 28858
rect 72114 28806 72166 28858
rect 67548 28704 67600 28756
rect 64880 28636 64932 28688
rect 67364 28636 67416 28688
rect 67548 28568 67600 28620
rect 67364 28500 67416 28552
rect 74210 28262 74262 28314
rect 74274 28262 74326 28314
rect 74338 28262 74390 28314
rect 74402 28262 74454 28314
rect 74466 28262 74518 28314
rect 65892 27820 65944 27872
rect 63500 27732 63552 27784
rect 71858 27718 71910 27770
rect 71922 27718 71974 27770
rect 71986 27718 72038 27770
rect 72050 27718 72102 27770
rect 72114 27718 72166 27770
rect 68192 27548 68244 27600
rect 67548 27412 67600 27464
rect 74210 27174 74262 27226
rect 74274 27174 74326 27226
rect 74338 27174 74390 27226
rect 74402 27174 74454 27226
rect 74466 27174 74518 27226
rect 64880 27072 64932 27124
rect 68100 27072 68152 27124
rect 66628 27047 66680 27056
rect 66628 27013 66637 27047
rect 66637 27013 66671 27047
rect 66671 27013 66680 27047
rect 66628 27004 66680 27013
rect 70676 26936 70728 26988
rect 71858 26630 71910 26682
rect 71922 26630 71974 26682
rect 71986 26630 72038 26682
rect 72050 26630 72102 26682
rect 72114 26630 72166 26682
rect 63500 26528 63552 26580
rect 67640 26528 67692 26580
rect 67364 26324 67416 26376
rect 63408 26256 63460 26308
rect 63500 26188 63552 26240
rect 63408 26052 63460 26104
rect 74210 26086 74262 26138
rect 74274 26086 74326 26138
rect 74338 26086 74390 26138
rect 74402 26086 74454 26138
rect 74466 26086 74518 26138
rect 63592 25984 63644 26036
rect 63500 25780 63552 25832
rect 63592 25780 63644 25832
rect 63684 25712 63736 25764
rect 65432 25644 65484 25696
rect 71858 25542 71910 25594
rect 71922 25542 71974 25594
rect 71986 25542 72038 25594
rect 72050 25542 72102 25594
rect 72114 25542 72166 25594
rect 68652 25440 68704 25492
rect 74210 24998 74262 25050
rect 74274 24998 74326 25050
rect 74338 24998 74390 25050
rect 74402 24998 74454 25050
rect 74466 24998 74518 25050
rect 71858 24454 71910 24506
rect 71922 24454 71974 24506
rect 71986 24454 72038 24506
rect 72050 24454 72102 24506
rect 72114 24454 72166 24506
rect 67732 24352 67784 24404
rect 65156 24284 65208 24336
rect 66444 24148 66496 24200
rect 74210 23910 74262 23962
rect 74274 23910 74326 23962
rect 74338 23910 74390 23962
rect 74402 23910 74454 23962
rect 74466 23910 74518 23962
rect 64972 23808 65024 23860
rect 67640 23604 67692 23656
rect 65524 23468 65576 23520
rect 71858 23366 71910 23418
rect 71922 23366 71974 23418
rect 71986 23366 72038 23418
rect 72050 23366 72102 23418
rect 72114 23366 72166 23418
rect 68284 23264 68336 23316
rect 68836 23196 68888 23248
rect 66444 23060 66496 23112
rect 74210 22822 74262 22874
rect 74274 22822 74326 22874
rect 74338 22822 74390 22874
rect 74402 22822 74454 22874
rect 74466 22822 74518 22874
rect 71858 22278 71910 22330
rect 71922 22278 71974 22330
rect 71986 22278 72038 22330
rect 72050 22278 72102 22330
rect 72114 22278 72166 22330
rect 66444 22176 66496 22228
rect 67732 22176 67784 22228
rect 65156 22108 65208 22160
rect 74210 21734 74262 21786
rect 74274 21734 74326 21786
rect 74338 21734 74390 21786
rect 74402 21734 74454 21786
rect 74466 21734 74518 21786
rect 69388 21496 69440 21548
rect 71858 21190 71910 21242
rect 71922 21190 71974 21242
rect 71986 21190 72038 21242
rect 72050 21190 72102 21242
rect 72114 21190 72166 21242
rect 68192 21088 68244 21140
rect 74210 20646 74262 20698
rect 74274 20646 74326 20698
rect 74338 20646 74390 20698
rect 74402 20646 74454 20698
rect 74466 20646 74518 20698
rect 65156 20204 65208 20256
rect 71858 20102 71910 20154
rect 71922 20102 71974 20154
rect 71986 20102 72038 20154
rect 72050 20102 72102 20154
rect 72114 20102 72166 20154
rect 74210 19558 74262 19610
rect 74274 19558 74326 19610
rect 74338 19558 74390 19610
rect 74402 19558 74454 19610
rect 74466 19558 74518 19610
rect 65064 19116 65116 19168
rect 71858 19014 71910 19066
rect 71922 19014 71974 19066
rect 71986 19014 72038 19066
rect 72050 19014 72102 19066
rect 72114 19014 72166 19066
rect 67824 18912 67876 18964
rect 74210 18470 74262 18522
rect 74274 18470 74326 18522
rect 74338 18470 74390 18522
rect 74402 18470 74454 18522
rect 74466 18470 74518 18522
rect 65156 17960 65208 18012
rect 71858 17926 71910 17978
rect 71922 17926 71974 17978
rect 71986 17926 72038 17978
rect 72050 17926 72102 17978
rect 72114 17926 72166 17978
rect 74210 17382 74262 17434
rect 74274 17382 74326 17434
rect 74338 17382 74390 17434
rect 74402 17382 74454 17434
rect 74466 17382 74518 17434
rect 65616 16940 65668 16992
rect 71858 16838 71910 16890
rect 71922 16838 71974 16890
rect 71986 16838 72038 16890
rect 72050 16838 72102 16890
rect 72114 16838 72166 16890
rect 63408 16600 63460 16652
rect 63408 16396 63460 16448
rect 63776 16396 63828 16448
rect 74210 16294 74262 16346
rect 74274 16294 74326 16346
rect 74338 16294 74390 16346
rect 74402 16294 74454 16346
rect 74466 16294 74518 16346
rect 71858 15750 71910 15802
rect 71922 15750 71974 15802
rect 71986 15750 72038 15802
rect 72050 15750 72102 15802
rect 72114 15750 72166 15802
rect 65156 15580 65208 15632
rect 74210 15206 74262 15258
rect 74274 15206 74326 15258
rect 74338 15206 74390 15258
rect 74402 15206 74454 15258
rect 74466 15206 74518 15258
rect 64972 14764 65024 14816
rect 71858 14662 71910 14714
rect 71922 14662 71974 14714
rect 71986 14662 72038 14714
rect 72050 14662 72102 14714
rect 72114 14662 72166 14714
rect 67640 14560 67692 14612
rect 74210 14118 74262 14170
rect 74274 14118 74326 14170
rect 74338 14118 74390 14170
rect 74402 14118 74454 14170
rect 74466 14118 74518 14170
rect 65156 13676 65208 13728
rect 71858 13574 71910 13626
rect 71922 13574 71974 13626
rect 71986 13574 72038 13626
rect 72050 13574 72102 13626
rect 72114 13574 72166 13626
rect 74210 13030 74262 13082
rect 74274 13030 74326 13082
rect 74338 13030 74390 13082
rect 74402 13030 74454 13082
rect 74466 13030 74518 13082
rect 64880 12724 64932 12776
rect 67732 12588 67784 12640
rect 71858 12486 71910 12538
rect 71922 12486 71974 12538
rect 71986 12486 72038 12538
rect 72050 12486 72102 12538
rect 72114 12486 72166 12538
rect 63408 12112 63460 12164
rect 63868 12112 63920 12164
rect 74210 11942 74262 11994
rect 74274 11942 74326 11994
rect 74338 11942 74390 11994
rect 74402 11942 74454 11994
rect 74466 11942 74518 11994
rect 63500 11840 63552 11892
rect 63776 11840 63828 11892
rect 71858 11398 71910 11450
rect 71922 11398 71974 11450
rect 71986 11398 72038 11450
rect 72050 11398 72102 11450
rect 72114 11398 72166 11450
rect 65156 11228 65208 11280
rect 64052 11024 64104 11076
rect 66812 11024 66864 11076
rect 74210 10854 74262 10906
rect 74274 10854 74326 10906
rect 74338 10854 74390 10906
rect 74402 10854 74454 10906
rect 74466 10854 74518 10906
rect 64880 10412 64932 10464
rect 63408 10292 63460 10344
rect 71858 10310 71910 10362
rect 71922 10310 71974 10362
rect 71986 10310 72038 10362
rect 72050 10310 72102 10362
rect 72114 10310 72166 10362
rect 74210 9766 74262 9818
rect 74274 9766 74326 9818
rect 74338 9766 74390 9818
rect 74402 9766 74454 9818
rect 74466 9766 74518 9818
rect 65156 9324 65208 9376
rect 71858 9222 71910 9274
rect 71922 9222 71974 9274
rect 71986 9222 72038 9274
rect 72050 9222 72102 9274
rect 72114 9222 72166 9274
rect 74210 8678 74262 8730
rect 74274 8678 74326 8730
rect 74338 8678 74390 8730
rect 74402 8678 74454 8730
rect 74466 8678 74518 8730
rect 71858 8134 71910 8186
rect 71922 8134 71974 8186
rect 71986 8134 72038 8186
rect 72050 8134 72102 8186
rect 72114 8134 72166 8186
rect 62948 7828 63000 7880
rect 65616 7828 65668 7880
rect 52276 7760 52328 7812
rect 60740 7760 60792 7812
rect 61660 7760 61712 7812
rect 64604 7760 64656 7812
rect 43536 7692 43588 7744
rect 62764 7692 62816 7744
rect 62856 7692 62908 7744
rect 64972 7692 65024 7744
rect 48044 7624 48096 7676
rect 24584 7556 24636 7608
rect 55588 7624 55640 7676
rect 63408 7624 63460 7676
rect 54852 7556 54904 7608
rect 65064 7556 65116 7608
rect 74210 7590 74262 7642
rect 74274 7590 74326 7642
rect 74338 7590 74390 7642
rect 74402 7590 74454 7642
rect 74466 7590 74518 7642
rect 54668 7420 54720 7472
rect 60740 7488 60792 7540
rect 67824 7488 67876 7540
rect 62764 7420 62816 7472
rect 68100 7420 68152 7472
rect 63500 7352 63552 7404
rect 60740 7284 60792 7336
rect 65708 7284 65760 7336
rect 62672 7216 62724 7268
rect 65800 7216 65852 7268
rect 59084 7148 59136 7200
rect 65892 7148 65944 7200
rect 60464 7080 60516 7132
rect 64604 7080 64656 7132
rect 55772 6944 55824 6996
rect 65064 7012 65116 7064
rect 71858 7046 71910 7098
rect 71922 7046 71974 7098
rect 71986 7046 72038 7098
rect 72050 7046 72102 7098
rect 72114 7046 72166 7098
rect 54668 6876 54720 6928
rect 46112 6808 46164 6860
rect 55864 6808 55916 6860
rect 61016 6876 61068 6928
rect 60556 6808 60608 6860
rect 61384 6808 61436 6860
rect 64880 6808 64932 6860
rect 65800 6808 65852 6860
rect 66720 6808 66772 6860
rect 69388 6808 69440 6860
rect 48872 6740 48924 6792
rect 63684 6740 63736 6792
rect 64972 6740 65024 6792
rect 67916 6740 67968 6792
rect 42616 6672 42668 6724
rect 27528 6604 27580 6656
rect 61384 6604 61436 6656
rect 23296 6536 23348 6588
rect 62948 6536 63000 6588
rect 65708 6672 65760 6724
rect 67088 6672 67140 6724
rect 65064 6604 65116 6656
rect 68836 6604 68888 6656
rect 64972 6536 65024 6588
rect 28908 6468 28960 6520
rect 46388 6468 46440 6520
rect 51724 6468 51776 6520
rect 55772 6468 55824 6520
rect 55864 6468 55916 6520
rect 64696 6468 64748 6520
rect 74210 6502 74262 6554
rect 74274 6502 74326 6554
rect 74338 6502 74390 6554
rect 74402 6502 74454 6554
rect 74466 6502 74518 6554
rect 24768 6400 24820 6452
rect 60832 6400 60884 6452
rect 61016 6400 61068 6452
rect 63408 6400 63460 6452
rect 63684 6400 63736 6452
rect 66260 6400 66312 6452
rect 32956 6332 33008 6384
rect 48228 6332 48280 6384
rect 54852 6332 54904 6384
rect 67732 6332 67784 6384
rect 23664 6264 23716 6316
rect 32864 6264 32916 6316
rect 51080 6264 51132 6316
rect 63960 6264 64012 6316
rect 64972 6264 65024 6316
rect 68652 6264 68704 6316
rect 27068 6196 27120 6248
rect 45652 6196 45704 6248
rect 48136 6196 48188 6248
rect 24952 6128 25004 6180
rect 44916 6128 44968 6180
rect 47032 6128 47084 6180
rect 51080 6128 51132 6180
rect 53288 6196 53340 6248
rect 57428 6196 57480 6248
rect 57520 6196 57572 6248
rect 60464 6196 60516 6248
rect 60648 6196 60700 6248
rect 63868 6196 63920 6248
rect 64696 6196 64748 6248
rect 66996 6196 67048 6248
rect 63776 6128 63828 6180
rect 64604 6128 64656 6180
rect 68376 6128 68428 6180
rect 26148 6060 26200 6112
rect 34888 6060 34940 6112
rect 45560 6060 45612 6112
rect 55680 6060 55732 6112
rect 55864 6060 55916 6112
rect 62856 6060 62908 6112
rect 63408 6060 63460 6112
rect 68192 6060 68244 6112
rect 1858 5958 1910 6010
rect 1922 5958 1974 6010
rect 1986 5958 2038 6010
rect 2050 5958 2102 6010
rect 2114 5958 2166 6010
rect 11858 5958 11910 6010
rect 11922 5958 11974 6010
rect 11986 5958 12038 6010
rect 12050 5958 12102 6010
rect 12114 5958 12166 6010
rect 21858 5958 21910 6010
rect 21922 5958 21974 6010
rect 21986 5958 22038 6010
rect 22050 5958 22102 6010
rect 22114 5958 22166 6010
rect 31858 5958 31910 6010
rect 31922 5958 31974 6010
rect 31986 5958 32038 6010
rect 32050 5958 32102 6010
rect 32114 5958 32166 6010
rect 41858 5958 41910 6010
rect 41922 5958 41974 6010
rect 41986 5958 42038 6010
rect 42050 5958 42102 6010
rect 42114 5958 42166 6010
rect 51858 5958 51910 6010
rect 51922 5958 51974 6010
rect 51986 5958 52038 6010
rect 52050 5958 52102 6010
rect 52114 5958 52166 6010
rect 61858 5958 61910 6010
rect 61922 5958 61974 6010
rect 61986 5958 62038 6010
rect 62050 5958 62102 6010
rect 62114 5958 62166 6010
rect 71858 5958 71910 6010
rect 71922 5958 71974 6010
rect 71986 5958 72038 6010
rect 72050 5958 72102 6010
rect 72114 5958 72166 6010
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 26148 5899 26200 5908
rect 26148 5865 26157 5899
rect 26157 5865 26191 5899
rect 26191 5865 26200 5899
rect 26148 5856 26200 5865
rect 29552 5856 29604 5908
rect 47492 5856 47544 5908
rect 48136 5899 48188 5908
rect 48136 5865 48145 5899
rect 48145 5865 48179 5899
rect 48179 5865 48188 5899
rect 48136 5856 48188 5865
rect 48872 5899 48924 5908
rect 48872 5865 48881 5899
rect 48881 5865 48915 5899
rect 48915 5865 48924 5899
rect 48872 5856 48924 5865
rect 53288 5856 53340 5908
rect 55864 5788 55916 5840
rect 57428 5856 57480 5908
rect 60832 5856 60884 5908
rect 62580 5856 62632 5908
rect 62764 5856 62816 5908
rect 63408 5856 63460 5908
rect 63776 5856 63828 5908
rect 65248 5856 65300 5908
rect 24584 5720 24636 5772
rect 24768 5763 24820 5772
rect 24768 5729 24777 5763
rect 24777 5729 24811 5763
rect 24811 5729 24820 5763
rect 24768 5720 24820 5729
rect 25044 5720 25096 5772
rect 32220 5720 32272 5772
rect 33876 5720 33928 5772
rect 25596 5652 25648 5704
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 25964 5695 26016 5704
rect 25964 5661 25973 5695
rect 25973 5661 26007 5695
rect 26007 5661 26016 5695
rect 25964 5652 26016 5661
rect 40408 5695 40460 5704
rect 40408 5661 40417 5695
rect 40417 5661 40451 5695
rect 40451 5661 40460 5695
rect 40408 5652 40460 5661
rect 41604 5652 41656 5704
rect 43536 5695 43588 5704
rect 43536 5661 43545 5695
rect 43545 5661 43579 5695
rect 43579 5661 43588 5695
rect 43536 5652 43588 5661
rect 43628 5652 43680 5704
rect 44640 5652 44692 5704
rect 44916 5763 44968 5772
rect 44916 5729 44925 5763
rect 44925 5729 44959 5763
rect 44959 5729 44968 5763
rect 44916 5720 44968 5729
rect 49792 5720 49844 5772
rect 51724 5720 51776 5772
rect 55220 5763 55272 5772
rect 55220 5729 55229 5763
rect 55229 5729 55263 5763
rect 55263 5729 55272 5763
rect 55220 5720 55272 5729
rect 56508 5763 56560 5772
rect 56508 5729 56517 5763
rect 56517 5729 56551 5763
rect 56551 5729 56560 5763
rect 56508 5720 56560 5729
rect 57796 5763 57848 5772
rect 57796 5729 57805 5763
rect 57805 5729 57839 5763
rect 57839 5729 57848 5763
rect 57796 5720 57848 5729
rect 58164 5763 58216 5772
rect 58164 5729 58173 5763
rect 58173 5729 58207 5763
rect 58207 5729 58216 5763
rect 58164 5720 58216 5729
rect 59452 5720 59504 5772
rect 45560 5695 45612 5704
rect 45560 5661 45569 5695
rect 45569 5661 45603 5695
rect 45603 5661 45612 5695
rect 45560 5652 45612 5661
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 46388 5695 46440 5704
rect 46388 5661 46397 5695
rect 46397 5661 46431 5695
rect 46431 5661 46440 5695
rect 46388 5652 46440 5661
rect 47032 5695 47084 5704
rect 47032 5661 47041 5695
rect 47041 5661 47075 5695
rect 47075 5661 47084 5695
rect 47032 5652 47084 5661
rect 47492 5695 47544 5704
rect 47492 5661 47501 5695
rect 47501 5661 47535 5695
rect 47535 5661 47544 5695
rect 47492 5652 47544 5661
rect 48228 5695 48280 5704
rect 48228 5661 48237 5695
rect 48237 5661 48271 5695
rect 48271 5661 48280 5695
rect 48228 5652 48280 5661
rect 50436 5695 50488 5704
rect 50436 5661 50445 5695
rect 50445 5661 50479 5695
rect 50479 5661 50488 5695
rect 50436 5652 50488 5661
rect 51264 5695 51316 5704
rect 51264 5661 51273 5695
rect 51273 5661 51307 5695
rect 51307 5661 51316 5695
rect 51264 5652 51316 5661
rect 52276 5652 52328 5704
rect 25044 5516 25096 5568
rect 31576 5516 31628 5568
rect 37004 5627 37056 5636
rect 37004 5593 37013 5627
rect 37013 5593 37047 5627
rect 37047 5593 37056 5627
rect 37004 5584 37056 5593
rect 49516 5584 49568 5636
rect 52368 5584 52420 5636
rect 33324 5516 33376 5568
rect 35900 5516 35952 5568
rect 41696 5559 41748 5568
rect 41696 5525 41705 5559
rect 41705 5525 41739 5559
rect 41739 5525 41748 5559
rect 41696 5516 41748 5525
rect 45928 5516 45980 5568
rect 47400 5516 47452 5568
rect 52552 5516 52604 5568
rect 52920 5652 52972 5704
rect 53840 5652 53892 5704
rect 56416 5652 56468 5704
rect 60740 5652 60792 5704
rect 61660 5763 61712 5772
rect 61660 5729 61669 5763
rect 61669 5729 61703 5763
rect 61703 5729 61712 5763
rect 61660 5720 61712 5729
rect 62580 5720 62632 5772
rect 67640 5788 67692 5840
rect 65984 5720 66036 5772
rect 66168 5763 66220 5772
rect 66168 5729 66177 5763
rect 66177 5729 66211 5763
rect 66211 5729 66220 5763
rect 66168 5720 66220 5729
rect 68468 5763 68520 5772
rect 68468 5729 68477 5763
rect 68477 5729 68511 5763
rect 68511 5729 68520 5763
rect 68468 5720 68520 5729
rect 53012 5584 53064 5636
rect 60924 5584 60976 5636
rect 61108 5584 61160 5636
rect 54668 5516 54720 5568
rect 54852 5516 54904 5568
rect 55588 5516 55640 5568
rect 56232 5516 56284 5568
rect 56324 5516 56376 5568
rect 59636 5516 59688 5568
rect 61200 5516 61252 5568
rect 62948 5695 63000 5704
rect 62948 5661 62957 5695
rect 62957 5661 62991 5695
rect 62991 5661 63000 5695
rect 62948 5652 63000 5661
rect 63592 5584 63644 5636
rect 65340 5584 65392 5636
rect 63316 5559 63368 5568
rect 63316 5525 63325 5559
rect 63325 5525 63359 5559
rect 63359 5525 63368 5559
rect 63316 5516 63368 5525
rect 64788 5516 64840 5568
rect 66444 5516 66496 5568
rect 68100 5559 68152 5568
rect 68100 5525 68109 5559
rect 68109 5525 68143 5559
rect 68143 5525 68152 5559
rect 68100 5516 68152 5525
rect 4210 5414 4262 5466
rect 4274 5414 4326 5466
rect 4338 5414 4390 5466
rect 4402 5414 4454 5466
rect 4466 5414 4518 5466
rect 14210 5414 14262 5466
rect 14274 5414 14326 5466
rect 14338 5414 14390 5466
rect 14402 5414 14454 5466
rect 14466 5414 14518 5466
rect 24210 5414 24262 5466
rect 24274 5414 24326 5466
rect 24338 5414 24390 5466
rect 24402 5414 24454 5466
rect 24466 5414 24518 5466
rect 34210 5414 34262 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 44210 5414 44262 5466
rect 44274 5414 44326 5466
rect 44338 5414 44390 5466
rect 44402 5414 44454 5466
rect 44466 5414 44518 5466
rect 54210 5414 54262 5466
rect 54274 5414 54326 5466
rect 54338 5414 54390 5466
rect 54402 5414 54454 5466
rect 54466 5414 54518 5466
rect 64210 5414 64262 5466
rect 64274 5414 64326 5466
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 74210 5414 74262 5466
rect 74274 5414 74326 5466
rect 74338 5414 74390 5466
rect 74402 5414 74454 5466
rect 74466 5414 74518 5466
rect 26608 5312 26660 5364
rect 63592 5312 63644 5364
rect 23940 5176 23992 5228
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 25596 5219 25648 5228
rect 25596 5185 25605 5219
rect 25605 5185 25639 5219
rect 25639 5185 25648 5219
rect 25596 5176 25648 5185
rect 25964 5176 26016 5228
rect 26792 5244 26844 5296
rect 31208 5244 31260 5296
rect 24584 5108 24636 5160
rect 25412 5151 25464 5160
rect 25412 5117 25421 5151
rect 25421 5117 25455 5151
rect 25455 5117 25464 5151
rect 25412 5108 25464 5117
rect 25872 5151 25924 5160
rect 25872 5117 25881 5151
rect 25881 5117 25915 5151
rect 25915 5117 25924 5151
rect 25872 5108 25924 5117
rect 26608 5108 26660 5160
rect 23480 5040 23532 5092
rect 26792 5040 26844 5092
rect 27528 5151 27580 5160
rect 27528 5117 27537 5151
rect 27537 5117 27571 5151
rect 27571 5117 27580 5151
rect 27528 5108 27580 5117
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 28172 5176 28224 5228
rect 27988 5108 28040 5160
rect 28448 5219 28500 5228
rect 28448 5185 28457 5219
rect 28457 5185 28491 5219
rect 28491 5185 28500 5219
rect 28448 5176 28500 5185
rect 29644 5219 29696 5228
rect 29644 5185 29653 5219
rect 29653 5185 29687 5219
rect 29687 5185 29696 5219
rect 29644 5176 29696 5185
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 29000 5040 29052 5092
rect 30288 5151 30340 5160
rect 30288 5117 30297 5151
rect 30297 5117 30331 5151
rect 30331 5117 30340 5151
rect 30288 5108 30340 5117
rect 30380 5108 30432 5160
rect 46204 5244 46256 5296
rect 46480 5244 46532 5296
rect 59084 5244 59136 5296
rect 61016 5244 61068 5296
rect 62856 5244 62908 5296
rect 69664 5244 69716 5296
rect 31392 5176 31444 5228
rect 40408 5151 40460 5160
rect 40408 5117 40417 5151
rect 40417 5117 40451 5151
rect 40451 5117 40460 5151
rect 40408 5108 40460 5117
rect 41052 5151 41104 5160
rect 41052 5117 41061 5151
rect 41061 5117 41095 5151
rect 41095 5117 41104 5151
rect 41052 5108 41104 5117
rect 41512 5151 41564 5160
rect 41512 5117 41521 5151
rect 41521 5117 41555 5151
rect 41555 5117 41564 5151
rect 41512 5108 41564 5117
rect 42984 5219 43036 5228
rect 42984 5185 42993 5219
rect 42993 5185 43027 5219
rect 43027 5185 43036 5219
rect 42984 5176 43036 5185
rect 45928 5176 45980 5228
rect 46296 5219 46348 5228
rect 46296 5185 46305 5219
rect 46305 5185 46339 5219
rect 46339 5185 46348 5219
rect 46296 5176 46348 5185
rect 44088 5108 44140 5160
rect 44640 5108 44692 5160
rect 45376 5151 45428 5160
rect 45376 5117 45385 5151
rect 45385 5117 45419 5151
rect 45419 5117 45428 5151
rect 45376 5108 45428 5117
rect 46020 5108 46072 5160
rect 46388 5108 46440 5160
rect 47492 5151 47544 5160
rect 47492 5117 47501 5151
rect 47501 5117 47535 5151
rect 47535 5117 47544 5151
rect 47492 5108 47544 5117
rect 48044 5108 48096 5160
rect 49148 5151 49200 5160
rect 49148 5117 49157 5151
rect 49157 5117 49191 5151
rect 49191 5117 49200 5151
rect 49148 5108 49200 5117
rect 49792 5151 49844 5160
rect 49792 5117 49801 5151
rect 49801 5117 49835 5151
rect 49835 5117 49844 5151
rect 49792 5108 49844 5117
rect 52368 5176 52420 5228
rect 53012 5176 53064 5228
rect 53104 5219 53156 5228
rect 53104 5185 53113 5219
rect 53113 5185 53147 5219
rect 53147 5185 53156 5219
rect 53104 5176 53156 5185
rect 54576 5176 54628 5228
rect 53288 5151 53340 5160
rect 53288 5117 53297 5151
rect 53297 5117 53331 5151
rect 53331 5117 53340 5151
rect 53288 5108 53340 5117
rect 53380 5108 53432 5160
rect 54944 5219 54996 5228
rect 54944 5185 54953 5219
rect 54953 5185 54987 5219
rect 54987 5185 54996 5219
rect 54944 5176 54996 5185
rect 55036 5176 55088 5228
rect 56416 5108 56468 5160
rect 61292 5176 61344 5228
rect 65432 5108 65484 5160
rect 69940 5108 69992 5160
rect 29276 5040 29328 5092
rect 29644 5040 29696 5092
rect 26148 4972 26200 5024
rect 26240 5015 26292 5024
rect 26240 4981 26249 5015
rect 26249 4981 26283 5015
rect 26283 4981 26292 5015
rect 26240 4972 26292 4981
rect 26700 5015 26752 5024
rect 26700 4981 26709 5015
rect 26709 4981 26743 5015
rect 26743 4981 26752 5015
rect 26700 4972 26752 4981
rect 27804 4972 27856 5024
rect 27896 5015 27948 5024
rect 27896 4981 27905 5015
rect 27905 4981 27939 5015
rect 27939 4981 27948 5015
rect 27896 4972 27948 4981
rect 28540 4972 28592 5024
rect 28724 5015 28776 5024
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 28816 4972 28868 5024
rect 29092 4972 29144 5024
rect 29368 5015 29420 5024
rect 29368 4981 29377 5015
rect 29377 4981 29411 5015
rect 29411 4981 29420 5015
rect 29368 4972 29420 4981
rect 29460 4972 29512 5024
rect 30472 5015 30524 5024
rect 30472 4981 30481 5015
rect 30481 4981 30515 5015
rect 30515 4981 30524 5015
rect 30472 4972 30524 4981
rect 45008 4972 45060 5024
rect 45100 5015 45152 5024
rect 45100 4981 45109 5015
rect 45109 4981 45143 5015
rect 45143 4981 45152 5015
rect 45100 4972 45152 4981
rect 46112 4972 46164 5024
rect 47032 5040 47084 5092
rect 47308 5040 47360 5092
rect 63776 5040 63828 5092
rect 69756 5040 69808 5092
rect 47124 4972 47176 5024
rect 47400 4972 47452 5024
rect 49332 4972 49384 5024
rect 52920 5015 52972 5024
rect 52920 4981 52929 5015
rect 52929 4981 52963 5015
rect 52963 4981 52972 5015
rect 52920 4972 52972 4981
rect 54668 4972 54720 5024
rect 54760 4972 54812 5024
rect 63500 4972 63552 5024
rect 69848 4972 69900 5024
rect 71412 4972 71464 5024
rect 73252 5015 73304 5024
rect 73252 4981 73261 5015
rect 73261 4981 73295 5015
rect 73295 4981 73304 5015
rect 73252 4972 73304 4981
rect 1858 4870 1910 4922
rect 1922 4870 1974 4922
rect 1986 4870 2038 4922
rect 2050 4870 2102 4922
rect 2114 4870 2166 4922
rect 11858 4870 11910 4922
rect 11922 4870 11974 4922
rect 11986 4870 12038 4922
rect 12050 4870 12102 4922
rect 12114 4870 12166 4922
rect 21858 4870 21910 4922
rect 21922 4870 21974 4922
rect 21986 4870 22038 4922
rect 22050 4870 22102 4922
rect 22114 4870 22166 4922
rect 31858 4870 31910 4922
rect 31922 4870 31974 4922
rect 31986 4870 32038 4922
rect 32050 4870 32102 4922
rect 32114 4870 32166 4922
rect 41858 4870 41910 4922
rect 41922 4870 41974 4922
rect 41986 4870 42038 4922
rect 42050 4870 42102 4922
rect 42114 4870 42166 4922
rect 51858 4870 51910 4922
rect 51922 4870 51974 4922
rect 51986 4870 52038 4922
rect 52050 4870 52102 4922
rect 52114 4870 52166 4922
rect 61858 4870 61910 4922
rect 61922 4870 61974 4922
rect 61986 4870 62038 4922
rect 62050 4870 62102 4922
rect 62114 4870 62166 4922
rect 71858 4870 71910 4922
rect 71922 4870 71974 4922
rect 71986 4870 72038 4922
rect 72050 4870 72102 4922
rect 72114 4870 72166 4922
rect 26240 4768 26292 4820
rect 30012 4768 30064 4820
rect 32312 4768 32364 4820
rect 41512 4768 41564 4820
rect 42616 4811 42668 4820
rect 42616 4777 42625 4811
rect 42625 4777 42659 4811
rect 42659 4777 42668 4811
rect 42616 4768 42668 4777
rect 45100 4768 45152 4820
rect 61016 4768 61068 4820
rect 62764 4768 62816 4820
rect 68744 4768 68796 4820
rect 25596 4700 25648 4752
rect 27712 4700 27764 4752
rect 27896 4700 27948 4752
rect 24584 4632 24636 4684
rect 31392 4632 31444 4684
rect 34060 4632 34112 4684
rect 35072 4700 35124 4752
rect 42984 4700 43036 4752
rect 36820 4632 36872 4684
rect 44732 4700 44784 4752
rect 45008 4700 45060 4752
rect 26700 4564 26752 4616
rect 29000 4564 29052 4616
rect 29092 4564 29144 4616
rect 25412 4496 25464 4548
rect 30104 4496 30156 4548
rect 26148 4428 26200 4480
rect 29644 4428 29696 4480
rect 33968 4607 34020 4616
rect 33968 4573 33977 4607
rect 33977 4573 34011 4607
rect 34011 4573 34020 4607
rect 33968 4564 34020 4573
rect 41236 4607 41288 4616
rect 41236 4573 41245 4607
rect 41245 4573 41279 4607
rect 41279 4573 41288 4607
rect 41236 4564 41288 4573
rect 41696 4564 41748 4616
rect 43352 4607 43404 4616
rect 43352 4573 43361 4607
rect 43361 4573 43395 4607
rect 43395 4573 43404 4607
rect 43352 4564 43404 4573
rect 32588 4496 32640 4548
rect 36544 4496 36596 4548
rect 46296 4564 46348 4616
rect 46664 4607 46716 4616
rect 46664 4573 46673 4607
rect 46673 4573 46707 4607
rect 46707 4573 46716 4607
rect 46664 4564 46716 4573
rect 47032 4632 47084 4684
rect 49332 4700 49384 4752
rect 65156 4700 65208 4752
rect 34704 4428 34756 4480
rect 43904 4428 43956 4480
rect 46572 4496 46624 4548
rect 45928 4428 45980 4480
rect 46756 4428 46808 4480
rect 48964 4496 49016 4548
rect 51540 4632 51592 4684
rect 54852 4632 54904 4684
rect 54944 4632 54996 4684
rect 70768 4632 70820 4684
rect 61016 4564 61068 4616
rect 61292 4564 61344 4616
rect 61476 4564 61528 4616
rect 68560 4564 68612 4616
rect 60924 4496 60976 4548
rect 49056 4428 49108 4480
rect 55496 4428 55548 4480
rect 61108 4471 61160 4480
rect 61108 4437 61117 4471
rect 61117 4437 61151 4471
rect 61151 4437 61160 4471
rect 61108 4428 61160 4437
rect 62856 4496 62908 4548
rect 69296 4496 69348 4548
rect 68008 4428 68060 4480
rect 4210 4326 4262 4378
rect 4274 4326 4326 4378
rect 4338 4326 4390 4378
rect 4402 4326 4454 4378
rect 4466 4326 4518 4378
rect 14210 4326 14262 4378
rect 14274 4326 14326 4378
rect 14338 4326 14390 4378
rect 14402 4326 14454 4378
rect 14466 4326 14518 4378
rect 24210 4326 24262 4378
rect 24274 4326 24326 4378
rect 24338 4326 24390 4378
rect 24402 4326 24454 4378
rect 24466 4326 24518 4378
rect 34210 4326 34262 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 44210 4326 44262 4378
rect 44274 4326 44326 4378
rect 44338 4326 44390 4378
rect 44402 4326 44454 4378
rect 44466 4326 44518 4378
rect 54210 4326 54262 4378
rect 54274 4326 54326 4378
rect 54338 4326 54390 4378
rect 54402 4326 54454 4378
rect 54466 4326 54518 4378
rect 64210 4326 64262 4378
rect 64274 4326 64326 4378
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 74210 4326 74262 4378
rect 74274 4326 74326 4378
rect 74338 4326 74390 4378
rect 74402 4326 74454 4378
rect 74466 4326 74518 4378
rect 27620 4224 27672 4276
rect 34796 4224 34848 4276
rect 36544 4224 36596 4276
rect 47492 4224 47544 4276
rect 47584 4224 47636 4276
rect 51540 4224 51592 4276
rect 53288 4224 53340 4276
rect 62672 4224 62724 4276
rect 19064 4088 19116 4140
rect 20260 4088 20312 4140
rect 27620 4131 27672 4140
rect 27620 4097 27629 4131
rect 27629 4097 27663 4131
rect 27663 4097 27672 4131
rect 27620 4088 27672 4097
rect 30104 4156 30156 4208
rect 27988 4020 28040 4072
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 31484 4088 31536 4140
rect 34612 4088 34664 4140
rect 34704 4131 34756 4140
rect 34704 4097 34713 4131
rect 34713 4097 34747 4131
rect 34747 4097 34756 4131
rect 34704 4088 34756 4097
rect 34796 4088 34848 4140
rect 34980 4088 35032 4140
rect 42984 4088 43036 4140
rect 43904 4088 43956 4140
rect 47032 4088 47084 4140
rect 65524 4156 65576 4208
rect 48964 4088 49016 4140
rect 55496 4088 55548 4140
rect 60740 4088 60792 4140
rect 66628 4088 66680 4140
rect 41696 4020 41748 4072
rect 61476 4020 61528 4072
rect 66536 4020 66588 4072
rect 17868 3952 17920 4004
rect 40408 3952 40460 4004
rect 47032 3952 47084 4004
rect 51264 3952 51316 4004
rect 60924 3952 60976 4004
rect 62764 3952 62816 4004
rect 23388 3884 23440 3936
rect 27620 3884 27672 3936
rect 33968 3884 34020 3936
rect 34796 3884 34848 3936
rect 35808 3884 35860 3936
rect 37004 3884 37056 3936
rect 47400 3884 47452 3936
rect 1858 3782 1910 3834
rect 1922 3782 1974 3834
rect 1986 3782 2038 3834
rect 2050 3782 2102 3834
rect 2114 3782 2166 3834
rect 11858 3782 11910 3834
rect 11922 3782 11974 3834
rect 11986 3782 12038 3834
rect 12050 3782 12102 3834
rect 12114 3782 12166 3834
rect 21858 3782 21910 3834
rect 21922 3782 21974 3834
rect 21986 3782 22038 3834
rect 22050 3782 22102 3834
rect 22114 3782 22166 3834
rect 31858 3782 31910 3834
rect 31922 3782 31974 3834
rect 31986 3782 32038 3834
rect 32050 3782 32102 3834
rect 32114 3782 32166 3834
rect 41858 3782 41910 3834
rect 41922 3782 41974 3834
rect 41986 3782 42038 3834
rect 42050 3782 42102 3834
rect 42114 3782 42166 3834
rect 51858 3782 51910 3834
rect 51922 3782 51974 3834
rect 51986 3782 52038 3834
rect 52050 3782 52102 3834
rect 52114 3782 52166 3834
rect 61858 3782 61910 3834
rect 61922 3782 61974 3834
rect 61986 3782 62038 3834
rect 62050 3782 62102 3834
rect 62114 3782 62166 3834
rect 71858 3782 71910 3834
rect 71922 3782 71974 3834
rect 71986 3782 72038 3834
rect 72050 3782 72102 3834
rect 72114 3782 72166 3834
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20904 3680 20956 3732
rect 25596 3680 25648 3732
rect 26056 3723 26108 3732
rect 26056 3689 26065 3723
rect 26065 3689 26099 3723
rect 26099 3689 26108 3723
rect 26056 3680 26108 3689
rect 29736 3680 29788 3732
rect 25780 3612 25832 3664
rect 32312 3680 32364 3732
rect 32680 3612 32732 3664
rect 18236 3476 18288 3528
rect 20536 3476 20588 3528
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 22468 3476 22520 3528
rect 23388 3476 23440 3528
rect 24952 3519 25004 3528
rect 24952 3485 24961 3519
rect 24961 3485 24995 3519
rect 24995 3485 25004 3519
rect 24952 3476 25004 3485
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 25780 3519 25832 3528
rect 25780 3485 25789 3519
rect 25789 3485 25823 3519
rect 25823 3485 25832 3519
rect 25780 3476 25832 3485
rect 25964 3476 26016 3528
rect 27896 3544 27948 3596
rect 28172 3544 28224 3596
rect 32772 3544 32824 3596
rect 33232 3680 33284 3732
rect 41236 3680 41288 3732
rect 36176 3612 36228 3664
rect 49148 3612 49200 3664
rect 28724 3476 28776 3528
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31576 3476 31628 3528
rect 32220 3519 32272 3528
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 32864 3519 32916 3528
rect 32864 3485 32873 3519
rect 32873 3485 32907 3519
rect 32907 3485 32916 3519
rect 32864 3476 32916 3485
rect 36084 3544 36136 3596
rect 44640 3544 44692 3596
rect 20628 3340 20680 3392
rect 25596 3408 25648 3460
rect 27712 3451 27764 3460
rect 27712 3417 27721 3451
rect 27721 3417 27755 3451
rect 27755 3417 27764 3451
rect 27712 3408 27764 3417
rect 37096 3476 37148 3528
rect 42248 3476 42300 3528
rect 52552 3544 52604 3596
rect 55864 3544 55916 3596
rect 66352 3544 66404 3596
rect 51172 3476 51224 3528
rect 67364 3476 67416 3528
rect 23112 3340 23164 3392
rect 23296 3383 23348 3392
rect 23296 3349 23305 3383
rect 23305 3349 23339 3383
rect 23339 3349 23348 3383
rect 23296 3340 23348 3349
rect 26240 3340 26292 3392
rect 27160 3340 27212 3392
rect 45376 3408 45428 3460
rect 27896 3383 27948 3392
rect 27896 3349 27905 3383
rect 27905 3349 27939 3383
rect 27939 3349 27948 3383
rect 27896 3340 27948 3349
rect 27988 3340 28040 3392
rect 31300 3340 31352 3392
rect 31392 3383 31444 3392
rect 31392 3349 31401 3383
rect 31401 3349 31435 3383
rect 31435 3349 31444 3383
rect 31392 3340 31444 3349
rect 39764 3340 39816 3392
rect 44916 3340 44968 3392
rect 61384 3408 61436 3460
rect 4210 3238 4262 3290
rect 4274 3238 4326 3290
rect 4338 3238 4390 3290
rect 4402 3238 4454 3290
rect 4466 3238 4518 3290
rect 14210 3238 14262 3290
rect 14274 3238 14326 3290
rect 14338 3238 14390 3290
rect 14402 3238 14454 3290
rect 14466 3238 14518 3290
rect 24210 3238 24262 3290
rect 24274 3238 24326 3290
rect 24338 3238 24390 3290
rect 24402 3238 24454 3290
rect 24466 3238 24518 3290
rect 34210 3238 34262 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 44210 3238 44262 3290
rect 44274 3238 44326 3290
rect 44338 3238 44390 3290
rect 44402 3238 44454 3290
rect 44466 3238 44518 3290
rect 54210 3238 54262 3290
rect 54274 3238 54326 3290
rect 54338 3238 54390 3290
rect 54402 3238 54454 3290
rect 54466 3238 54518 3290
rect 64210 3238 64262 3290
rect 64274 3238 64326 3290
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 74210 3238 74262 3290
rect 74274 3238 74326 3290
rect 74338 3238 74390 3290
rect 74402 3238 74454 3290
rect 74466 3238 74518 3290
rect 20536 3179 20588 3188
rect 20536 3145 20545 3179
rect 20545 3145 20579 3179
rect 20579 3145 20588 3179
rect 20536 3136 20588 3145
rect 24860 3136 24912 3188
rect 25780 3136 25832 3188
rect 27712 3136 27764 3188
rect 29552 3136 29604 3188
rect 17868 3111 17920 3120
rect 17868 3077 17877 3111
rect 17877 3077 17911 3111
rect 17911 3077 17920 3111
rect 17868 3068 17920 3077
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 20720 3000 20772 3052
rect 18696 2932 18748 2984
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 22744 3000 22796 3052
rect 20536 2864 20588 2916
rect 21732 2975 21784 2984
rect 21732 2941 21741 2975
rect 21741 2941 21775 2975
rect 21775 2941 21784 2975
rect 21732 2932 21784 2941
rect 22284 2864 22336 2916
rect 22928 3068 22980 3120
rect 26056 3068 26108 3120
rect 23112 3043 23164 3052
rect 23112 3009 23121 3043
rect 23121 3009 23155 3043
rect 23155 3009 23164 3043
rect 23112 3000 23164 3009
rect 29368 3068 29420 3120
rect 33232 3136 33284 3188
rect 34980 3136 35032 3188
rect 36728 3136 36780 3188
rect 37004 3179 37056 3188
rect 37004 3145 37013 3179
rect 37013 3145 37047 3179
rect 37047 3145 37056 3179
rect 37004 3136 37056 3145
rect 37096 3068 37148 3120
rect 42432 3068 42484 3120
rect 64696 3068 64748 3120
rect 23020 2932 23072 2984
rect 24032 2932 24084 2984
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 26240 2864 26292 2916
rect 26976 3000 27028 3052
rect 27160 3000 27212 3052
rect 27068 2975 27120 2984
rect 27068 2941 27077 2975
rect 27077 2941 27111 2975
rect 27111 2941 27120 2975
rect 27068 2932 27120 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 28908 2975 28960 2984
rect 28908 2941 28917 2975
rect 28917 2941 28951 2975
rect 28951 2941 28960 2975
rect 28908 2932 28960 2941
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 29552 3043 29604 3052
rect 29552 3009 29561 3043
rect 29561 3009 29595 3043
rect 29595 3009 29604 3043
rect 29552 3000 29604 3009
rect 29644 3000 29696 3052
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 31484 3000 31536 3052
rect 31668 3000 31720 3052
rect 32312 3000 32364 3052
rect 33140 3000 33192 3052
rect 33324 3043 33376 3052
rect 33324 3009 33333 3043
rect 33333 3009 33367 3043
rect 33367 3009 33376 3043
rect 33324 3000 33376 3009
rect 30196 2932 30248 2984
rect 32220 2975 32272 2984
rect 32220 2941 32229 2975
rect 32229 2941 32263 2975
rect 32263 2941 32272 2975
rect 32220 2932 32272 2941
rect 29460 2864 29512 2916
rect 34060 3043 34112 3052
rect 34060 3009 34069 3043
rect 34069 3009 34103 3043
rect 34103 3009 34112 3043
rect 34060 3000 34112 3009
rect 34612 3000 34664 3052
rect 34888 3043 34940 3052
rect 34888 3009 34897 3043
rect 34897 3009 34931 3043
rect 34931 3009 34940 3043
rect 34888 3000 34940 3009
rect 36176 3000 36228 3052
rect 36636 3000 36688 3052
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 34796 2932 34848 2984
rect 35808 2975 35860 2984
rect 35808 2941 35817 2975
rect 35817 2941 35851 2975
rect 35851 2941 35860 2975
rect 35808 2932 35860 2941
rect 37096 2932 37148 2984
rect 45928 3043 45980 3052
rect 45928 3009 45937 3043
rect 45937 3009 45971 3043
rect 45971 3009 45980 3043
rect 45928 3000 45980 3009
rect 47124 3000 47176 3052
rect 49056 3043 49108 3052
rect 49056 3009 49065 3043
rect 49065 3009 49099 3043
rect 49099 3009 49108 3043
rect 49056 3000 49108 3009
rect 52920 3043 52972 3052
rect 52920 3009 52929 3043
rect 52929 3009 52963 3043
rect 52963 3009 52972 3043
rect 52920 3000 52972 3009
rect 53932 3000 53984 3052
rect 54668 3043 54720 3052
rect 54668 3009 54677 3043
rect 54677 3009 54711 3043
rect 54711 3009 54720 3043
rect 54668 3000 54720 3009
rect 56232 3043 56284 3052
rect 56232 3009 56241 3043
rect 56241 3009 56275 3043
rect 56275 3009 56284 3043
rect 56232 3000 56284 3009
rect 57796 3043 57848 3052
rect 57796 3009 57805 3043
rect 57805 3009 57839 3043
rect 57839 3009 57848 3043
rect 57796 3000 57848 3009
rect 59452 3043 59504 3052
rect 59452 3009 59461 3043
rect 59461 3009 59495 3043
rect 59495 3009 59504 3043
rect 59452 3000 59504 3009
rect 61200 3043 61252 3052
rect 61200 3009 61209 3043
rect 61209 3009 61243 3043
rect 61243 3009 61252 3043
rect 61200 3000 61252 3009
rect 63224 3043 63276 3052
rect 63224 3009 63233 3043
rect 63233 3009 63267 3043
rect 63267 3009 63276 3043
rect 63224 3000 63276 3009
rect 64788 3043 64840 3052
rect 64788 3009 64797 3043
rect 64797 3009 64831 3043
rect 64831 3009 64840 3043
rect 64788 3000 64840 3009
rect 66444 3043 66496 3052
rect 66444 3009 66453 3043
rect 66453 3009 66487 3043
rect 66487 3009 66496 3043
rect 66444 3000 66496 3009
rect 68100 3043 68152 3052
rect 68100 3009 68109 3043
rect 68109 3009 68143 3043
rect 68143 3009 68152 3043
rect 68100 3000 68152 3009
rect 69848 3043 69900 3052
rect 69848 3009 69857 3043
rect 69857 3009 69891 3043
rect 69891 3009 69900 3043
rect 69848 3000 69900 3009
rect 71412 3043 71464 3052
rect 71412 3009 71421 3043
rect 71421 3009 71455 3043
rect 71455 3009 71464 3043
rect 71412 3000 71464 3009
rect 73252 3000 73304 3052
rect 63592 2932 63644 2984
rect 44824 2864 44876 2916
rect 50068 2864 50120 2916
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 22560 2796 22612 2848
rect 24952 2839 25004 2848
rect 24952 2805 24961 2839
rect 24961 2805 24995 2839
rect 24995 2805 25004 2839
rect 24952 2796 25004 2805
rect 25964 2839 26016 2848
rect 25964 2805 25973 2839
rect 25973 2805 26007 2839
rect 26007 2805 26016 2839
rect 25964 2796 26016 2805
rect 26516 2839 26568 2848
rect 26516 2805 26525 2839
rect 26525 2805 26559 2839
rect 26559 2805 26568 2839
rect 26516 2796 26568 2805
rect 28172 2796 28224 2848
rect 30932 2839 30984 2848
rect 30932 2805 30941 2839
rect 30941 2805 30975 2839
rect 30975 2805 30984 2839
rect 30932 2796 30984 2805
rect 32588 2796 32640 2848
rect 32956 2796 33008 2848
rect 33876 2796 33928 2848
rect 34704 2796 34756 2848
rect 35808 2796 35860 2848
rect 44916 2796 44968 2848
rect 47584 2796 47636 2848
rect 52644 2796 52696 2848
rect 53104 2839 53156 2848
rect 53104 2805 53113 2839
rect 53113 2805 53147 2839
rect 53147 2805 53156 2839
rect 53104 2796 53156 2805
rect 55220 2796 55272 2848
rect 56416 2839 56468 2848
rect 56416 2805 56425 2839
rect 56425 2805 56459 2839
rect 56459 2805 56468 2839
rect 56416 2796 56468 2805
rect 57980 2839 58032 2848
rect 57980 2805 57989 2839
rect 57989 2805 58023 2839
rect 58023 2805 58032 2839
rect 57980 2796 58032 2805
rect 60372 2796 60424 2848
rect 61384 2839 61436 2848
rect 61384 2805 61393 2839
rect 61393 2805 61427 2839
rect 61427 2805 61436 2839
rect 61384 2796 61436 2805
rect 63040 2839 63092 2848
rect 63040 2805 63049 2839
rect 63049 2805 63083 2839
rect 63083 2805 63092 2839
rect 63040 2796 63092 2805
rect 64604 2839 64656 2848
rect 64604 2805 64613 2839
rect 64613 2805 64647 2839
rect 64647 2805 64656 2839
rect 64604 2796 64656 2805
rect 66260 2839 66312 2848
rect 66260 2805 66269 2839
rect 66269 2805 66303 2839
rect 66303 2805 66312 2839
rect 66260 2796 66312 2805
rect 68284 2839 68336 2848
rect 68284 2805 68293 2839
rect 68293 2805 68327 2839
rect 68327 2805 68336 2839
rect 68284 2796 68336 2805
rect 69664 2839 69716 2848
rect 69664 2805 69673 2839
rect 69673 2805 69707 2839
rect 69707 2805 69716 2839
rect 69664 2796 69716 2805
rect 71228 2839 71280 2848
rect 71228 2805 71237 2839
rect 71237 2805 71271 2839
rect 71271 2805 71280 2839
rect 71228 2796 71280 2805
rect 73252 2796 73304 2848
rect 1858 2694 1910 2746
rect 1922 2694 1974 2746
rect 1986 2694 2038 2746
rect 2050 2694 2102 2746
rect 2114 2694 2166 2746
rect 11858 2694 11910 2746
rect 11922 2694 11974 2746
rect 11986 2694 12038 2746
rect 12050 2694 12102 2746
rect 12114 2694 12166 2746
rect 21858 2694 21910 2746
rect 21922 2694 21974 2746
rect 21986 2694 22038 2746
rect 22050 2694 22102 2746
rect 22114 2694 22166 2746
rect 31858 2694 31910 2746
rect 31922 2694 31974 2746
rect 31986 2694 32038 2746
rect 32050 2694 32102 2746
rect 32114 2694 32166 2746
rect 41858 2694 41910 2746
rect 41922 2694 41974 2746
rect 41986 2694 42038 2746
rect 42050 2694 42102 2746
rect 42114 2694 42166 2746
rect 51858 2694 51910 2746
rect 51922 2694 51974 2746
rect 51986 2694 52038 2746
rect 52050 2694 52102 2746
rect 52114 2694 52166 2746
rect 61858 2694 61910 2746
rect 61922 2694 61974 2746
rect 61986 2694 62038 2746
rect 62050 2694 62102 2746
rect 62114 2694 62166 2746
rect 71858 2694 71910 2746
rect 71922 2694 71974 2746
rect 71986 2694 72038 2746
rect 72050 2694 72102 2746
rect 72114 2694 72166 2746
rect 18144 2592 18196 2644
rect 19156 2592 19208 2644
rect 19892 2635 19944 2644
rect 19892 2601 19901 2635
rect 19901 2601 19935 2635
rect 19935 2601 19944 2635
rect 19892 2592 19944 2601
rect 20812 2592 20864 2644
rect 21732 2592 21784 2644
rect 24032 2592 24084 2644
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 25320 2635 25372 2644
rect 25320 2601 25329 2635
rect 25329 2601 25363 2635
rect 25363 2601 25372 2635
rect 25320 2592 25372 2601
rect 27528 2635 27580 2644
rect 27528 2601 27537 2635
rect 27537 2601 27571 2635
rect 27571 2601 27580 2635
rect 27528 2592 27580 2601
rect 29092 2592 29144 2644
rect 16948 2388 17000 2440
rect 23296 2524 23348 2576
rect 25872 2524 25924 2576
rect 30472 2524 30524 2576
rect 19708 2456 19760 2508
rect 20812 2456 20864 2508
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 20168 2388 20220 2440
rect 20536 2320 20588 2372
rect 21364 2388 21416 2440
rect 25964 2456 26016 2508
rect 27804 2456 27856 2508
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 24032 2388 24084 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2388 25280 2440
rect 26056 2431 26108 2440
rect 26056 2397 26065 2431
rect 26065 2397 26099 2431
rect 26099 2397 26108 2431
rect 26056 2388 26108 2397
rect 26148 2388 26200 2440
rect 26884 2388 26936 2440
rect 27436 2388 27488 2440
rect 28448 2456 28500 2508
rect 70676 2592 70728 2644
rect 31668 2567 31720 2576
rect 31668 2533 31677 2567
rect 31677 2533 31711 2567
rect 31711 2533 31720 2567
rect 31668 2524 31720 2533
rect 33140 2567 33192 2576
rect 33140 2533 33149 2567
rect 33149 2533 33183 2567
rect 33183 2533 33192 2567
rect 33140 2524 33192 2533
rect 34060 2524 34112 2576
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 35440 2456 35492 2508
rect 39396 2524 39448 2576
rect 43352 2524 43404 2576
rect 44732 2524 44784 2576
rect 51172 2524 51224 2576
rect 53932 2567 53984 2576
rect 53932 2533 53941 2567
rect 53941 2533 53975 2567
rect 53975 2533 53984 2567
rect 53932 2524 53984 2533
rect 54024 2524 54076 2576
rect 28632 2431 28684 2440
rect 28632 2397 28641 2431
rect 28641 2397 28675 2431
rect 28675 2397 28684 2431
rect 28632 2388 28684 2397
rect 29184 2388 29236 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 32220 2388 32272 2440
rect 32496 2431 32548 2440
rect 32496 2397 32505 2431
rect 32505 2397 32539 2431
rect 32539 2397 32548 2431
rect 32496 2388 32548 2397
rect 33600 2431 33652 2440
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 47860 2456 47912 2508
rect 48044 2456 48096 2508
rect 55312 2456 55364 2508
rect 41696 2388 41748 2440
rect 42340 2388 42392 2440
rect 43444 2388 43496 2440
rect 45560 2431 45612 2440
rect 45560 2397 45569 2431
rect 45569 2397 45603 2431
rect 45603 2397 45612 2431
rect 45560 2388 45612 2397
rect 46204 2431 46256 2440
rect 46204 2397 46213 2431
rect 46213 2397 46247 2431
rect 46247 2397 46256 2431
rect 46204 2388 46256 2397
rect 47308 2388 47360 2440
rect 21732 2320 21784 2372
rect 17776 2252 17828 2304
rect 17868 2252 17920 2304
rect 20904 2252 20956 2304
rect 26700 2295 26752 2304
rect 26700 2261 26709 2295
rect 26709 2261 26743 2295
rect 26743 2261 26752 2295
rect 26700 2252 26752 2261
rect 28540 2295 28592 2304
rect 28540 2261 28549 2295
rect 28549 2261 28583 2295
rect 28583 2261 28592 2295
rect 28540 2252 28592 2261
rect 29092 2252 29144 2304
rect 30288 2295 30340 2304
rect 30288 2261 30297 2295
rect 30297 2261 30331 2295
rect 30331 2261 30340 2295
rect 30288 2252 30340 2261
rect 31300 2252 31352 2304
rect 33048 2252 33100 2304
rect 35072 2252 35124 2304
rect 39120 2320 39172 2372
rect 43076 2363 43128 2372
rect 43076 2329 43085 2363
rect 43085 2329 43119 2363
rect 43119 2329 43128 2363
rect 43076 2320 43128 2329
rect 39396 2252 39448 2304
rect 39580 2252 39632 2304
rect 46388 2320 46440 2372
rect 46848 2252 46900 2304
rect 47216 2363 47268 2372
rect 47216 2329 47225 2363
rect 47225 2329 47259 2363
rect 47259 2329 47268 2363
rect 47216 2320 47268 2329
rect 49056 2431 49108 2440
rect 49056 2397 49065 2431
rect 49065 2397 49099 2431
rect 49099 2397 49108 2431
rect 49056 2388 49108 2397
rect 53840 2388 53892 2440
rect 53932 2388 53984 2440
rect 57336 2431 57388 2440
rect 57336 2397 57345 2431
rect 57345 2397 57379 2431
rect 57379 2397 57388 2431
rect 57336 2388 57388 2397
rect 53748 2320 53800 2372
rect 55036 2320 55088 2372
rect 56692 2320 56744 2372
rect 66168 2524 66220 2576
rect 65708 2456 65760 2508
rect 67456 2499 67508 2508
rect 67456 2465 67465 2499
rect 67465 2465 67499 2499
rect 67499 2465 67508 2499
rect 67456 2456 67508 2465
rect 49424 2252 49476 2304
rect 49516 2252 49568 2304
rect 54760 2295 54812 2304
rect 54760 2261 54769 2295
rect 54769 2261 54803 2295
rect 54803 2261 54812 2295
rect 54760 2252 54812 2261
rect 57888 2252 57940 2304
rect 60740 2320 60792 2372
rect 61016 2363 61068 2372
rect 61016 2329 61025 2363
rect 61025 2329 61059 2363
rect 61059 2329 61068 2363
rect 61016 2320 61068 2329
rect 62304 2431 62356 2440
rect 62304 2397 62313 2431
rect 62313 2397 62347 2431
rect 62347 2397 62356 2431
rect 62304 2388 62356 2397
rect 62948 2295 63000 2304
rect 62948 2261 62957 2295
rect 62957 2261 62991 2295
rect 62991 2261 63000 2295
rect 62948 2252 63000 2261
rect 63592 2320 63644 2372
rect 65524 2388 65576 2440
rect 67272 2388 67324 2440
rect 69940 2431 69992 2440
rect 69940 2397 69949 2431
rect 69949 2397 69983 2431
rect 69983 2397 69992 2431
rect 69940 2388 69992 2397
rect 70492 2388 70544 2440
rect 67548 2320 67600 2372
rect 63684 2252 63736 2304
rect 66076 2252 66128 2304
rect 69388 2252 69440 2304
rect 71044 2252 71096 2304
rect 4210 2150 4262 2202
rect 4274 2150 4326 2202
rect 4338 2150 4390 2202
rect 4402 2150 4454 2202
rect 4466 2150 4518 2202
rect 14210 2150 14262 2202
rect 14274 2150 14326 2202
rect 14338 2150 14390 2202
rect 14402 2150 14454 2202
rect 14466 2150 14518 2202
rect 24210 2150 24262 2202
rect 24274 2150 24326 2202
rect 24338 2150 24390 2202
rect 24402 2150 24454 2202
rect 24466 2150 24518 2202
rect 34210 2150 34262 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 44210 2150 44262 2202
rect 44274 2150 44326 2202
rect 44338 2150 44390 2202
rect 44402 2150 44454 2202
rect 44466 2150 44518 2202
rect 54210 2150 54262 2202
rect 54274 2150 54326 2202
rect 54338 2150 54390 2202
rect 54402 2150 54454 2202
rect 54466 2150 54518 2202
rect 64210 2150 64262 2202
rect 64274 2150 64326 2202
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 74210 2150 74262 2202
rect 74274 2150 74326 2202
rect 74338 2150 74390 2202
rect 74402 2150 74454 2202
rect 74466 2150 74518 2202
rect 17592 2048 17644 2100
rect 18236 2048 18288 2100
rect 17868 1980 17920 2032
rect 21456 2048 21508 2100
rect 24584 2048 24636 2100
rect 16396 1912 16448 1964
rect 18420 1912 18472 1964
rect 20260 1955 20312 1964
rect 20260 1921 20269 1955
rect 20269 1921 20303 1955
rect 20303 1921 20312 1955
rect 20260 1912 20312 1921
rect 21456 1955 21508 1964
rect 21456 1921 21465 1955
rect 21465 1921 21499 1955
rect 21499 1921 21508 1955
rect 21456 1912 21508 1921
rect 18052 1844 18104 1896
rect 22376 1912 22428 1964
rect 23480 1912 23532 1964
rect 24952 1912 25004 1964
rect 25872 1955 25924 1964
rect 25872 1921 25881 1955
rect 25881 1921 25915 1955
rect 25915 1921 25924 1955
rect 25872 1912 25924 1921
rect 26148 1955 26200 1964
rect 26148 1921 26157 1955
rect 26157 1921 26191 1955
rect 26191 1921 26200 1955
rect 26148 1912 26200 1921
rect 26700 1912 26752 1964
rect 28540 1980 28592 2032
rect 32312 2048 32364 2100
rect 32496 2091 32548 2100
rect 32496 2057 32505 2091
rect 32505 2057 32539 2091
rect 32539 2057 32548 2091
rect 32496 2048 32548 2057
rect 34612 2091 34664 2100
rect 34612 2057 34621 2091
rect 34621 2057 34655 2091
rect 34655 2057 34664 2091
rect 34612 2048 34664 2057
rect 36636 2048 36688 2100
rect 39120 2091 39172 2100
rect 39120 2057 39129 2091
rect 39129 2057 39163 2091
rect 39163 2057 39172 2091
rect 39120 2048 39172 2057
rect 41696 2048 41748 2100
rect 47032 2048 47084 2100
rect 48044 2048 48096 2100
rect 54024 2048 54076 2100
rect 55036 2091 55088 2100
rect 55036 2057 55045 2091
rect 55045 2057 55079 2091
rect 55079 2057 55088 2091
rect 55036 2048 55088 2057
rect 61476 2048 61528 2100
rect 63592 2091 63644 2100
rect 63592 2057 63601 2091
rect 63601 2057 63635 2091
rect 63635 2057 63644 2091
rect 63592 2048 63644 2057
rect 22836 1887 22888 1896
rect 22836 1853 22845 1887
rect 22845 1853 22879 1887
rect 22879 1853 22888 1887
rect 22836 1844 22888 1853
rect 24676 1844 24728 1896
rect 28448 1844 28500 1896
rect 21456 1776 21508 1828
rect 20628 1708 20680 1760
rect 26976 1708 27028 1760
rect 29092 1955 29144 1964
rect 29092 1921 29101 1955
rect 29101 1921 29135 1955
rect 29135 1921 29144 1955
rect 29092 1912 29144 1921
rect 29552 1912 29604 1964
rect 66904 1980 66956 2032
rect 67272 2091 67324 2100
rect 67272 2057 67281 2091
rect 67281 2057 67315 2091
rect 67315 2057 67324 2091
rect 67272 2048 67324 2057
rect 70584 2048 70636 2100
rect 69204 1980 69256 2032
rect 70124 1980 70176 2032
rect 29920 1912 29972 1964
rect 30288 1844 30340 1896
rect 31300 1955 31352 1964
rect 31300 1921 31309 1955
rect 31309 1921 31343 1955
rect 31343 1921 31352 1955
rect 31300 1912 31352 1921
rect 34060 1912 34112 1964
rect 34796 1955 34848 1964
rect 34796 1921 34805 1955
rect 34805 1921 34839 1955
rect 34839 1921 34848 1955
rect 34796 1912 34848 1921
rect 39028 1912 39080 1964
rect 42892 1912 42944 1964
rect 42984 1955 43036 1964
rect 42984 1921 42993 1955
rect 42993 1921 43027 1955
rect 43027 1921 43036 1955
rect 42984 1912 43036 1921
rect 32404 1844 32456 1896
rect 34612 1844 34664 1896
rect 36176 1887 36228 1896
rect 36176 1853 36185 1887
rect 36185 1853 36219 1887
rect 36219 1853 36228 1887
rect 36176 1844 36228 1853
rect 37556 1887 37608 1896
rect 37556 1853 37565 1887
rect 37565 1853 37599 1887
rect 37599 1853 37608 1887
rect 37556 1844 37608 1853
rect 41144 1887 41196 1896
rect 41144 1853 41153 1887
rect 41153 1853 41187 1887
rect 41187 1853 41196 1887
rect 41144 1844 41196 1853
rect 35900 1776 35952 1828
rect 42984 1776 43036 1828
rect 44916 1887 44968 1896
rect 44916 1853 44925 1887
rect 44925 1853 44959 1887
rect 44959 1853 44968 1887
rect 44916 1844 44968 1853
rect 45376 1955 45428 1964
rect 45376 1921 45385 1955
rect 45385 1921 45419 1955
rect 45419 1921 45428 1955
rect 45376 1912 45428 1921
rect 45652 1912 45704 1964
rect 46848 1912 46900 1964
rect 47584 1912 47636 1964
rect 49516 1955 49568 1964
rect 49516 1921 49525 1955
rect 49525 1921 49559 1955
rect 49559 1921 49568 1955
rect 49516 1912 49568 1921
rect 53104 1955 53156 1964
rect 53104 1921 53113 1955
rect 53113 1921 53147 1955
rect 53147 1921 53156 1955
rect 53104 1912 53156 1921
rect 54760 1912 54812 1964
rect 56416 1955 56468 1964
rect 56416 1921 56425 1955
rect 56425 1921 56459 1955
rect 56459 1921 56468 1955
rect 56416 1912 56468 1921
rect 57888 1955 57940 1964
rect 57888 1921 57897 1955
rect 57897 1921 57931 1955
rect 57931 1921 57940 1955
rect 57888 1912 57940 1921
rect 61384 1955 61436 1964
rect 61384 1921 61393 1955
rect 61393 1921 61427 1955
rect 61427 1921 61436 1955
rect 61384 1912 61436 1921
rect 62948 1955 63000 1964
rect 62948 1921 62957 1955
rect 62957 1921 62991 1955
rect 62991 1921 63000 1955
rect 62948 1912 63000 1921
rect 64604 1955 64656 1964
rect 64604 1921 64613 1955
rect 64613 1921 64647 1955
rect 64647 1921 64656 1955
rect 64604 1912 64656 1921
rect 66076 1955 66128 1964
rect 66076 1921 66085 1955
rect 66085 1921 66119 1955
rect 66119 1921 66128 1955
rect 66076 1912 66128 1921
rect 67180 1912 67232 1964
rect 69388 1955 69440 1964
rect 69388 1921 69397 1955
rect 69397 1921 69431 1955
rect 69431 1921 69440 1955
rect 69388 1912 69440 1921
rect 69664 1955 69716 1964
rect 69664 1921 69673 1955
rect 69673 1921 69707 1955
rect 69707 1921 69716 1955
rect 69664 1912 69716 1921
rect 71044 1955 71096 1964
rect 71044 1921 71053 1955
rect 71053 1921 71087 1955
rect 71087 1921 71096 1955
rect 71044 1912 71096 1921
rect 46020 1887 46072 1896
rect 46020 1853 46029 1887
rect 46029 1853 46063 1887
rect 46063 1853 46072 1887
rect 46020 1844 46072 1853
rect 46204 1887 46256 1896
rect 46204 1853 46213 1887
rect 46213 1853 46247 1887
rect 46247 1853 46256 1887
rect 46204 1844 46256 1853
rect 47860 1844 47912 1896
rect 51264 1887 51316 1896
rect 51264 1853 51273 1887
rect 51273 1853 51307 1887
rect 51307 1853 51316 1887
rect 51264 1844 51316 1853
rect 50436 1776 50488 1828
rect 39580 1708 39632 1760
rect 42248 1708 42300 1760
rect 52736 1776 52788 1828
rect 52920 1844 52972 1896
rect 55588 1887 55640 1896
rect 55588 1853 55597 1887
rect 55597 1853 55631 1887
rect 55631 1853 55640 1887
rect 55588 1844 55640 1853
rect 56140 1844 56192 1896
rect 59360 1844 59412 1896
rect 60556 1887 60608 1896
rect 60556 1853 60565 1887
rect 60565 1853 60599 1887
rect 60599 1853 60608 1887
rect 60556 1844 60608 1853
rect 61108 1844 61160 1896
rect 63868 1887 63920 1896
rect 63868 1853 63877 1887
rect 63877 1853 63911 1887
rect 63911 1853 63920 1887
rect 63868 1844 63920 1853
rect 64696 1844 64748 1896
rect 72240 1844 72292 1896
rect 55864 1776 55916 1828
rect 65800 1776 65852 1828
rect 69388 1776 69440 1828
rect 57244 1708 57296 1760
rect 62396 1708 62448 1760
rect 65156 1708 65208 1760
rect 73160 1708 73212 1760
rect 1858 1606 1910 1658
rect 1922 1606 1974 1658
rect 1986 1606 2038 1658
rect 2050 1606 2102 1658
rect 2114 1606 2166 1658
rect 11858 1606 11910 1658
rect 11922 1606 11974 1658
rect 11986 1606 12038 1658
rect 12050 1606 12102 1658
rect 12114 1606 12166 1658
rect 21858 1606 21910 1658
rect 21922 1606 21974 1658
rect 21986 1606 22038 1658
rect 22050 1606 22102 1658
rect 22114 1606 22166 1658
rect 31858 1606 31910 1658
rect 31922 1606 31974 1658
rect 31986 1606 32038 1658
rect 32050 1606 32102 1658
rect 32114 1606 32166 1658
rect 41858 1606 41910 1658
rect 41922 1606 41974 1658
rect 41986 1606 42038 1658
rect 42050 1606 42102 1658
rect 42114 1606 42166 1658
rect 51858 1606 51910 1658
rect 51922 1606 51974 1658
rect 51986 1606 52038 1658
rect 52050 1606 52102 1658
rect 52114 1606 52166 1658
rect 61858 1606 61910 1658
rect 61922 1606 61974 1658
rect 61986 1606 62038 1658
rect 62050 1606 62102 1658
rect 62114 1606 62166 1658
rect 71858 1606 71910 1658
rect 71922 1606 71974 1658
rect 71986 1606 72038 1658
rect 72050 1606 72102 1658
rect 72114 1606 72166 1658
rect 22928 1504 22980 1556
rect 26056 1504 26108 1556
rect 28632 1504 28684 1556
rect 31024 1504 31076 1556
rect 32680 1504 32732 1556
rect 37464 1504 37516 1556
rect 37556 1504 37608 1556
rect 41144 1504 41196 1556
rect 45376 1504 45428 1556
rect 45560 1504 45612 1556
rect 47216 1504 47268 1556
rect 51264 1504 51316 1556
rect 61016 1504 61068 1556
rect 63868 1504 63920 1556
rect 69940 1504 69992 1556
rect 19156 1368 19208 1420
rect 20260 1368 20312 1420
rect 31116 1436 31168 1488
rect 31300 1436 31352 1488
rect 41604 1436 41656 1488
rect 22836 1368 22888 1420
rect 5080 1343 5132 1352
rect 5080 1309 5089 1343
rect 5089 1309 5123 1343
rect 5123 1309 5132 1343
rect 5080 1300 5132 1309
rect 15292 1300 15344 1352
rect 17500 1300 17552 1352
rect 17776 1343 17828 1352
rect 17776 1309 17785 1343
rect 17785 1309 17819 1343
rect 17819 1309 17828 1343
rect 17776 1300 17828 1309
rect 3148 1232 3200 1284
rect 15844 1232 15896 1284
rect 15568 1207 15620 1216
rect 15568 1173 15577 1207
rect 15577 1173 15611 1207
rect 15611 1173 15620 1207
rect 15568 1164 15620 1173
rect 19064 1300 19116 1352
rect 19432 1275 19484 1284
rect 19432 1241 19441 1275
rect 19441 1241 19475 1275
rect 19475 1241 19484 1275
rect 19432 1232 19484 1241
rect 19800 1343 19852 1352
rect 19800 1309 19809 1343
rect 19809 1309 19843 1343
rect 19843 1309 19852 1343
rect 19800 1300 19852 1309
rect 22560 1300 22612 1352
rect 22284 1232 22336 1284
rect 23572 1232 23624 1284
rect 26332 1300 26384 1352
rect 25780 1275 25832 1284
rect 25780 1241 25789 1275
rect 25789 1241 25823 1275
rect 25823 1241 25832 1275
rect 25780 1232 25832 1241
rect 26516 1164 26568 1216
rect 27988 1368 28040 1420
rect 27804 1300 27856 1352
rect 28080 1300 28132 1352
rect 33048 1368 33100 1420
rect 29000 1300 29052 1352
rect 30380 1300 30432 1352
rect 33232 1343 33284 1352
rect 33232 1309 33241 1343
rect 33241 1309 33275 1343
rect 33275 1309 33284 1343
rect 33232 1300 33284 1309
rect 37924 1368 37976 1420
rect 41236 1368 41288 1420
rect 43076 1368 43128 1420
rect 33508 1300 33560 1352
rect 27896 1164 27948 1216
rect 31300 1232 31352 1284
rect 33140 1232 33192 1284
rect 33600 1164 33652 1216
rect 35624 1343 35676 1352
rect 35624 1309 35633 1343
rect 35633 1309 35667 1343
rect 35667 1309 35676 1343
rect 35624 1300 35676 1309
rect 37372 1343 37424 1352
rect 37372 1309 37381 1343
rect 37381 1309 37415 1343
rect 37415 1309 37424 1343
rect 37372 1300 37424 1309
rect 37464 1300 37516 1352
rect 39764 1343 39816 1352
rect 39764 1309 39773 1343
rect 39773 1309 39807 1343
rect 39807 1309 39816 1343
rect 39764 1300 39816 1309
rect 40776 1300 40828 1352
rect 42432 1343 42484 1352
rect 42432 1309 42441 1343
rect 42441 1309 42475 1343
rect 42475 1309 42484 1343
rect 42432 1300 42484 1309
rect 42892 1300 42944 1352
rect 44824 1368 44876 1420
rect 46204 1368 46256 1420
rect 49608 1368 49660 1420
rect 59452 1368 59504 1420
rect 62764 1368 62816 1420
rect 67732 1368 67784 1420
rect 71044 1368 71096 1420
rect 44732 1300 44784 1352
rect 44916 1343 44968 1352
rect 44916 1309 44925 1343
rect 44925 1309 44959 1343
rect 44959 1309 44968 1343
rect 44916 1300 44968 1309
rect 36176 1232 36228 1284
rect 36268 1232 36320 1284
rect 39580 1232 39632 1284
rect 43996 1232 44048 1284
rect 45100 1232 45152 1284
rect 47400 1300 47452 1352
rect 49424 1300 49476 1352
rect 50068 1343 50120 1352
rect 50068 1309 50077 1343
rect 50077 1309 50111 1343
rect 50111 1309 50120 1343
rect 50068 1300 50120 1309
rect 50620 1300 50672 1352
rect 52644 1343 52696 1352
rect 52644 1309 52653 1343
rect 52653 1309 52687 1343
rect 52687 1309 52696 1343
rect 52644 1300 52696 1309
rect 53840 1300 53892 1352
rect 51172 1232 51224 1284
rect 35716 1164 35768 1216
rect 46020 1164 46072 1216
rect 52276 1164 52328 1216
rect 55220 1343 55272 1352
rect 55220 1309 55229 1343
rect 55229 1309 55263 1343
rect 55263 1309 55272 1343
rect 55220 1300 55272 1309
rect 56692 1343 56744 1352
rect 56692 1309 56701 1343
rect 56701 1309 56735 1343
rect 56735 1309 56744 1343
rect 56692 1300 56744 1309
rect 57244 1343 57296 1352
rect 57244 1309 57253 1343
rect 57253 1309 57287 1343
rect 57287 1309 57296 1343
rect 57244 1300 57296 1309
rect 57980 1343 58032 1352
rect 57980 1309 57989 1343
rect 57989 1309 58023 1343
rect 58023 1309 58032 1343
rect 57980 1300 58032 1309
rect 59360 1343 59412 1352
rect 59360 1309 59369 1343
rect 59369 1309 59403 1343
rect 59403 1309 59412 1343
rect 59360 1300 59412 1309
rect 54576 1232 54628 1284
rect 57796 1232 57848 1284
rect 58900 1232 58952 1284
rect 60372 1343 60424 1352
rect 60372 1309 60381 1343
rect 60381 1309 60415 1343
rect 60415 1309 60424 1343
rect 60372 1300 60424 1309
rect 62396 1343 62448 1352
rect 62396 1309 62405 1343
rect 62405 1309 62439 1343
rect 62439 1309 62448 1343
rect 62396 1300 62448 1309
rect 63040 1343 63092 1352
rect 63040 1309 63049 1343
rect 63049 1309 63083 1343
rect 63083 1309 63092 1343
rect 63040 1300 63092 1309
rect 63868 1300 63920 1352
rect 65156 1300 65208 1352
rect 66260 1343 66312 1352
rect 66260 1309 66269 1343
rect 66269 1309 66303 1343
rect 66303 1309 66312 1343
rect 66260 1300 66312 1309
rect 68284 1343 68336 1352
rect 68284 1309 68293 1343
rect 68293 1309 68327 1343
rect 68327 1309 68336 1343
rect 68284 1300 68336 1309
rect 68836 1300 68888 1352
rect 71228 1343 71280 1352
rect 71228 1309 71237 1343
rect 71237 1309 71271 1343
rect 71271 1309 71280 1343
rect 71228 1300 71280 1309
rect 73160 1300 73212 1352
rect 73252 1343 73304 1352
rect 73252 1309 73261 1343
rect 73261 1309 73295 1343
rect 73295 1309 73304 1343
rect 73252 1300 73304 1309
rect 66076 1232 66128 1284
rect 70032 1232 70084 1284
rect 67364 1164 67416 1216
rect 72700 1164 72752 1216
rect 4210 1062 4262 1114
rect 4274 1062 4326 1114
rect 4338 1062 4390 1114
rect 4402 1062 4454 1114
rect 4466 1062 4518 1114
rect 14210 1062 14262 1114
rect 14274 1062 14326 1114
rect 14338 1062 14390 1114
rect 14402 1062 14454 1114
rect 14466 1062 14518 1114
rect 24210 1062 24262 1114
rect 24274 1062 24326 1114
rect 24338 1062 24390 1114
rect 24402 1062 24454 1114
rect 24466 1062 24518 1114
rect 34210 1062 34262 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 44210 1062 44262 1114
rect 44274 1062 44326 1114
rect 44338 1062 44390 1114
rect 44402 1062 44454 1114
rect 44466 1062 44518 1114
rect 54210 1062 54262 1114
rect 54274 1062 54326 1114
rect 54338 1062 54390 1114
rect 54402 1062 54454 1114
rect 54466 1062 54518 1114
rect 64210 1062 64262 1114
rect 64274 1062 64326 1114
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 74210 1062 74262 1114
rect 74274 1062 74326 1114
rect 74338 1062 74390 1114
rect 74402 1062 74454 1114
rect 74466 1062 74518 1114
rect 5080 960 5132 1012
rect 23940 960 23992 1012
rect 31392 960 31444 1012
rect 35624 960 35676 1012
rect 15568 892 15620 944
rect 20720 892 20772 944
rect 27804 892 27856 944
rect 28540 892 28592 944
rect 19432 824 19484 876
rect 43628 824 43680 876
<< metal2 >>
rect 64188 84588 64540 86000
rect 64188 84532 64216 84588
rect 64272 84532 64296 84588
rect 64352 84532 64376 84588
rect 64432 84532 64456 84588
rect 64512 84532 64540 84588
rect 64188 84508 64540 84532
rect 64188 84452 64216 84508
rect 64272 84452 64296 84508
rect 64352 84452 64376 84508
rect 64432 84452 64456 84508
rect 64512 84452 64540 84508
rect 64188 84428 64540 84452
rect 64188 84372 64216 84428
rect 64272 84372 64296 84428
rect 64352 84372 64376 84428
rect 64432 84372 64456 84428
rect 64512 84372 64540 84428
rect 64188 84348 64540 84372
rect 64188 84292 64216 84348
rect 64272 84292 64296 84348
rect 64352 84292 64376 84348
rect 64432 84292 64456 84348
rect 64512 84292 64540 84348
rect 64188 74588 64540 84292
rect 71836 85434 72188 86000
rect 71836 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 72188 85434
rect 71836 84346 72188 85382
rect 71836 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 72188 84346
rect 64880 84244 64932 84250
rect 64880 84186 64932 84192
rect 64892 81802 64920 84186
rect 71836 83258 72188 84294
rect 71836 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 72188 83258
rect 66996 83156 67048 83162
rect 66996 83098 67048 83104
rect 64880 81796 64932 81802
rect 64880 81738 64932 81744
rect 64892 79898 64920 81738
rect 64880 79892 64932 79898
rect 64880 79834 64932 79840
rect 64892 77722 64920 79834
rect 66444 78736 66496 78742
rect 66444 78678 66496 78684
rect 64880 77716 64932 77722
rect 64880 77658 64932 77664
rect 64892 75206 64920 77658
rect 66260 76560 66312 76566
rect 66260 76502 66312 76508
rect 64880 75200 64932 75206
rect 64880 75142 64932 75148
rect 64188 74532 64216 74588
rect 64272 74532 64296 74588
rect 64352 74532 64376 74588
rect 64432 74532 64456 74588
rect 64512 74532 64540 74588
rect 64188 74508 64540 74532
rect 64188 74452 64216 74508
rect 64272 74452 64296 74508
rect 64352 74452 64376 74508
rect 64432 74452 64456 74508
rect 64512 74452 64540 74508
rect 64188 74428 64540 74452
rect 64188 74372 64216 74428
rect 64272 74372 64296 74428
rect 64352 74372 64376 74428
rect 64432 74372 64456 74428
rect 64512 74372 64540 74428
rect 64188 74348 64540 74372
rect 64188 74292 64216 74348
rect 64272 74292 64296 74348
rect 64352 74292 64376 74348
rect 64432 74292 64456 74348
rect 64512 74292 64540 74348
rect 63684 69624 63736 69630
rect 63684 69566 63736 69572
rect 63592 60920 63644 60926
rect 63592 60862 63644 60868
rect 63500 52624 63552 52630
rect 63498 52592 63500 52601
rect 63552 52592 63554 52601
rect 63498 52527 63554 52536
rect 63500 50312 63552 50318
rect 63498 50280 63500 50289
rect 63552 50280 63554 50289
rect 63498 50215 63554 50224
rect 63408 48821 63460 48827
rect 63406 48784 63408 48793
rect 63460 48784 63462 48793
rect 63406 48719 63462 48728
rect 63500 48113 63552 48119
rect 63498 48104 63500 48113
rect 63552 48104 63554 48113
rect 63498 48039 63554 48048
rect 63500 32144 63552 32150
rect 63500 32086 63552 32092
rect 63512 27962 63540 32086
rect 63420 27934 63540 27962
rect 63420 26466 63448 27934
rect 63500 27784 63552 27790
rect 63500 27726 63552 27732
rect 63512 26586 63540 27726
rect 63500 26580 63552 26586
rect 63500 26522 63552 26528
rect 63420 26438 63540 26466
rect 63408 26308 63460 26314
rect 63408 26250 63460 26256
rect 63420 26110 63448 26250
rect 63512 26246 63540 26438
rect 63500 26240 63552 26246
rect 63500 26182 63552 26188
rect 63408 26104 63460 26110
rect 63408 26046 63460 26052
rect 63604 26042 63632 60862
rect 63696 26217 63724 69566
rect 64188 64588 64540 74292
rect 64892 73234 64920 75142
rect 66168 74112 66220 74118
rect 66168 74054 66220 74060
rect 64880 73228 64932 73234
rect 64880 73170 64932 73176
rect 64892 71126 64920 73170
rect 65984 71936 66036 71942
rect 65984 71878 66036 71884
rect 64880 71120 64932 71126
rect 64880 71062 64932 71068
rect 64892 69018 64920 71062
rect 65524 70032 65576 70038
rect 65524 69974 65576 69980
rect 64880 69012 64932 69018
rect 64880 68954 64932 68960
rect 64604 67652 64656 67658
rect 64604 67594 64656 67600
rect 64188 64532 64216 64588
rect 64272 64532 64296 64588
rect 64352 64532 64376 64588
rect 64432 64532 64456 64588
rect 64512 64532 64540 64588
rect 64188 64508 64540 64532
rect 64188 64452 64216 64508
rect 64272 64452 64296 64508
rect 64352 64452 64376 64508
rect 64432 64452 64456 64508
rect 64512 64452 64540 64508
rect 64188 64428 64540 64452
rect 64188 64372 64216 64428
rect 64272 64372 64296 64428
rect 64352 64372 64376 64428
rect 64432 64372 64456 64428
rect 64512 64372 64540 64428
rect 64188 64348 64540 64372
rect 64188 64292 64216 64348
rect 64272 64292 64296 64348
rect 64352 64292 64376 64348
rect 64432 64292 64456 64348
rect 64512 64292 64540 64348
rect 64188 54588 64540 64292
rect 64188 54532 64216 54588
rect 64272 54532 64296 54588
rect 64352 54532 64376 54588
rect 64432 54532 64456 54588
rect 64512 54532 64540 54588
rect 64188 54508 64540 54532
rect 64188 54452 64216 54508
rect 64272 54452 64296 54508
rect 64352 54452 64376 54508
rect 64432 54452 64456 54508
rect 64512 54452 64540 54508
rect 64188 54428 64540 54452
rect 64188 54372 64216 54428
rect 64272 54372 64296 54428
rect 64352 54372 64376 54428
rect 64432 54372 64456 54428
rect 64512 54372 64540 54428
rect 64188 54348 64540 54372
rect 64188 54292 64216 54348
rect 64272 54292 64296 54348
rect 64352 54292 64376 54348
rect 64432 54292 64456 54348
rect 64512 54292 64540 54348
rect 63868 47728 63920 47734
rect 63866 47696 63868 47705
rect 63920 47696 63922 47705
rect 63866 47631 63922 47640
rect 63960 45756 64012 45762
rect 63960 45698 64012 45704
rect 63868 45280 63920 45286
rect 63868 45222 63920 45228
rect 63776 29640 63828 29646
rect 63776 29582 63828 29588
rect 63682 26208 63738 26217
rect 63682 26143 63738 26152
rect 63592 26036 63644 26042
rect 63592 25978 63644 25984
rect 63500 25832 63552 25838
rect 63500 25774 63552 25780
rect 63592 25832 63644 25838
rect 63592 25774 63644 25780
rect 63408 16652 63460 16658
rect 63408 16594 63460 16600
rect 63420 16454 63448 16594
rect 63408 16448 63460 16454
rect 63408 16390 63460 16396
rect 63408 12164 63460 12170
rect 63408 12106 63460 12112
rect 63420 10713 63448 12106
rect 63512 11898 63540 25774
rect 63500 11892 63552 11898
rect 63500 11834 63552 11840
rect 63498 11792 63554 11801
rect 63498 11727 63554 11736
rect 63406 10704 63462 10713
rect 63406 10639 63462 10648
rect 63408 10344 63460 10350
rect 63408 10286 63460 10292
rect 1836 6010 2188 7944
rect 1836 5958 1858 6010
rect 1910 5958 1922 6010
rect 1974 5958 1986 6010
rect 2038 5958 2050 6010
rect 2102 5958 2114 6010
rect 2166 5958 2188 6010
rect 1836 4922 2188 5958
rect 1836 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 2188 4922
rect 1836 3834 2188 4870
rect 1836 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 2188 3834
rect 1836 2746 2188 3782
rect 1836 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 2188 2746
rect 1836 2236 2188 2694
rect 1836 2180 1864 2236
rect 1920 2180 1944 2236
rect 2000 2180 2024 2236
rect 2080 2180 2104 2236
rect 2160 2180 2188 2236
rect 1836 2156 2188 2180
rect 1836 2100 1864 2156
rect 1920 2100 1944 2156
rect 2000 2100 2024 2156
rect 2080 2100 2104 2156
rect 2160 2100 2188 2156
rect 1836 2076 2188 2100
rect 1836 2020 1864 2076
rect 1920 2020 1944 2076
rect 2000 2020 2024 2076
rect 2080 2020 2104 2076
rect 2160 2020 2188 2076
rect 1836 1996 2188 2020
rect 1836 1940 1864 1996
rect 1920 1940 1944 1996
rect 2000 1940 2024 1996
rect 2080 1940 2104 1996
rect 2160 1940 2188 1996
rect 1836 1658 2188 1940
rect 1836 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 2188 1658
rect 1836 1040 2188 1606
rect 4188 5466 4540 7944
rect 4188 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 4540 5466
rect 4188 4588 4540 5414
rect 4188 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4540 4588
rect 4188 4508 4540 4532
rect 4188 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4540 4508
rect 4188 4428 4540 4452
rect 4188 4378 4216 4428
rect 4272 4378 4296 4428
rect 4352 4378 4376 4428
rect 4432 4378 4456 4428
rect 4512 4378 4540 4428
rect 4188 4326 4210 4378
rect 4272 4372 4274 4378
rect 4454 4372 4456 4378
rect 4262 4348 4274 4372
rect 4326 4348 4338 4372
rect 4390 4348 4402 4372
rect 4454 4348 4466 4372
rect 4272 4326 4274 4348
rect 4454 4326 4456 4348
rect 4518 4326 4540 4378
rect 4188 4292 4216 4326
rect 4272 4292 4296 4326
rect 4352 4292 4376 4326
rect 4432 4292 4456 4326
rect 4512 4292 4540 4326
rect 4188 3290 4540 4292
rect 4188 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 4540 3290
rect 4188 2202 4540 3238
rect 4188 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 4540 2202
rect 3148 1284 3200 1290
rect 3148 1226 3200 1232
rect 3160 800 3188 1226
rect 4188 1114 4540 2150
rect 11836 6010 12188 7944
rect 11836 5958 11858 6010
rect 11910 5958 11922 6010
rect 11974 5958 11986 6010
rect 12038 5958 12050 6010
rect 12102 5958 12114 6010
rect 12166 5958 12188 6010
rect 11836 4922 12188 5958
rect 11836 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 12188 4922
rect 11836 3834 12188 4870
rect 11836 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 12188 3834
rect 11836 2746 12188 3782
rect 11836 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 12188 2746
rect 11836 2236 12188 2694
rect 11836 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 12188 2236
rect 11836 2156 12188 2180
rect 11836 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 12188 2156
rect 11836 2076 12188 2100
rect 11836 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 12188 2076
rect 11836 1996 12188 2020
rect 11836 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 12188 1996
rect 11836 1658 12188 1940
rect 11836 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 12188 1658
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 4188 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 4540 1114
rect 4188 1040 4540 1062
rect 5092 1018 5120 1294
rect 11836 1040 12188 1606
rect 14188 5466 14540 7944
rect 14188 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 14540 5466
rect 14188 4588 14540 5414
rect 14188 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 14540 4588
rect 14188 4508 14540 4532
rect 14188 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 14540 4508
rect 14188 4428 14540 4452
rect 14188 4378 14216 4428
rect 14272 4378 14296 4428
rect 14352 4378 14376 4428
rect 14432 4378 14456 4428
rect 14512 4378 14540 4428
rect 14188 4326 14210 4378
rect 14272 4372 14274 4378
rect 14454 4372 14456 4378
rect 14262 4348 14274 4372
rect 14326 4348 14338 4372
rect 14390 4348 14402 4372
rect 14454 4348 14466 4372
rect 14272 4326 14274 4348
rect 14454 4326 14456 4348
rect 14518 4326 14540 4378
rect 14188 4292 14216 4326
rect 14272 4292 14296 4326
rect 14352 4292 14376 4326
rect 14432 4292 14456 4326
rect 14512 4292 14540 4326
rect 14188 3290 14540 4292
rect 21836 6010 22188 7944
rect 23296 6588 23348 6594
rect 23296 6530 23348 6536
rect 21836 5958 21858 6010
rect 21910 5958 21922 6010
rect 21974 5958 21986 6010
rect 22038 5958 22050 6010
rect 22102 5958 22114 6010
rect 22166 5958 22188 6010
rect 21836 4922 22188 5958
rect 23308 5778 23336 6530
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 5914 23704 6258
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 24188 5466 24540 7944
rect 24584 7608 24636 7614
rect 24584 7550 24636 7556
rect 24596 5778 24624 7550
rect 30286 6896 30342 6905
rect 30286 6831 30342 6840
rect 29642 6760 29698 6769
rect 29642 6695 29698 6704
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 29274 6624 29330 6633
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24780 5778 24808 6394
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24188 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 24540 5466
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 21836 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 22188 4922
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 14738 3360 14794 3369
rect 14738 3295 14794 3304
rect 14188 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 14540 3290
rect 14188 2202 14540 3238
rect 14188 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 14540 2202
rect 14188 1114 14540 2150
rect 14188 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 14540 1114
rect 14188 1040 14540 1062
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 14752 800 14780 3295
rect 17880 3126 17908 3946
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 16396 1964 16448 1970
rect 16396 1906 16448 1912
rect 15292 1352 15344 1358
rect 15292 1294 15344 1300
rect 15304 800 15332 1294
rect 15844 1284 15896 1290
rect 15844 1226 15896 1232
rect 15568 1216 15620 1222
rect 15568 1158 15620 1164
rect 15580 950 15608 1158
rect 15568 944 15620 950
rect 15568 886 15620 892
rect 15856 800 15884 1226
rect 16408 800 16436 1906
rect 16960 800 16988 2382
rect 17604 2106 17632 2382
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17592 2100 17644 2106
rect 17592 2042 17644 2048
rect 17788 1358 17816 2246
rect 17880 2038 17908 2246
rect 18248 2106 18276 3470
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 18432 1970 18460 2790
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 17500 1352 17552 1358
rect 17500 1294 17552 1300
rect 17776 1352 17828 1358
rect 17776 1294 17828 1300
rect 17512 800 17540 1294
rect 18064 800 18092 1838
rect 18708 1442 18736 2926
rect 18616 1414 18736 1442
rect 18616 800 18644 1414
rect 19076 1358 19104 4082
rect 20272 3738 20300 4082
rect 21836 3834 22188 4870
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 21836 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 22188 3834
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20548 3194 20576 3470
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 3058 20668 3334
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19168 2650 19196 2926
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 19064 1352 19116 1358
rect 19064 1294 19116 1300
rect 19168 800 19196 1362
rect 19432 1284 19484 1290
rect 19432 1226 19484 1232
rect 19444 882 19472 1226
rect 19432 876 19484 882
rect 19432 818 19484 824
rect 19720 800 19748 2450
rect 19812 1358 19840 2790
rect 19904 2650 19932 2926
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 20180 1272 20208 2382
rect 20548 2378 20576 2858
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20272 1426 20300 1906
rect 20640 1766 20668 2994
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 20260 1420 20312 1426
rect 20260 1362 20312 1368
rect 20180 1244 20300 1272
rect 20272 800 20300 1244
rect 20732 950 20760 2994
rect 20824 2650 20852 3470
rect 20916 2990 20944 3674
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20720 944 20772 950
rect 20720 886 20772 892
rect 20824 800 20852 2450
rect 20916 2310 20944 2926
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21376 800 21404 2382
rect 21468 2106 21496 2790
rect 21744 2650 21772 2926
rect 21836 2746 22188 3782
rect 23400 3534 23428 3878
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 21836 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 22188 2746
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 21468 1834 21496 1906
rect 21456 1828 21508 1834
rect 21456 1770 21508 1776
rect 21744 898 21772 2314
rect 21836 2236 22188 2694
rect 21836 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 22188 2236
rect 21836 2156 22188 2180
rect 21836 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 22188 2156
rect 21836 2076 22188 2100
rect 21836 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 22188 2076
rect 21836 1996 22188 2020
rect 21836 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 22188 1996
rect 21836 1658 22188 1940
rect 21836 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 22188 1658
rect 21836 1040 22188 1606
rect 22296 1290 22324 2858
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22388 1970 22416 2790
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 22284 1284 22336 1290
rect 22284 1226 22336 1232
rect 21744 870 21956 898
rect 21928 800 21956 870
rect 22480 800 22508 3470
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 22928 3120 22980 3126
rect 22756 3068 22928 3074
rect 22756 3062 22980 3068
rect 22756 3058 22968 3062
rect 23124 3058 23152 3334
rect 22744 3052 22968 3058
rect 22796 3046 22968 3052
rect 23112 3052 23164 3058
rect 22744 2994 22796 3000
rect 23112 2994 23164 3000
rect 23020 2984 23072 2990
rect 23020 2926 23072 2932
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 1358 22600 2790
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 22848 1426 22876 1838
rect 22940 1562 22968 2382
rect 22928 1556 22980 1562
rect 22928 1498 22980 1504
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 23032 800 23060 2926
rect 23308 2582 23336 3334
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 23492 1970 23520 5034
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 23572 1284 23624 1290
rect 23572 1226 23624 1232
rect 23584 800 23612 1226
rect 23952 1018 23980 5170
rect 24188 4588 24540 5414
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24596 4690 24624 5102
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 24188 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 24540 4588
rect 24188 4508 24540 4532
rect 24188 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 24540 4508
rect 24188 4428 24540 4452
rect 24188 4378 24216 4428
rect 24272 4378 24296 4428
rect 24352 4378 24376 4428
rect 24432 4378 24456 4428
rect 24512 4378 24540 4428
rect 24188 4326 24210 4378
rect 24272 4372 24274 4378
rect 24454 4372 24456 4378
rect 24262 4348 24274 4372
rect 24326 4348 24338 4372
rect 24390 4348 24402 4372
rect 24454 4348 24466 4372
rect 24272 4326 24274 4348
rect 24454 4326 24456 4348
rect 24518 4326 24540 4378
rect 24188 4292 24216 4326
rect 24272 4292 24296 4326
rect 24352 4292 24376 4326
rect 24432 4292 24456 4326
rect 24512 4292 24540 4326
rect 24188 3290 24540 4292
rect 24188 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 24540 3290
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 24044 2650 24072 2926
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23940 1012 23992 1018
rect 23940 954 23992 960
rect 24044 898 24072 2382
rect 24188 2202 24540 3238
rect 24872 3194 24900 5170
rect 24964 3534 24992 6122
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 25870 5944 25926 5953
rect 26160 5914 26188 6054
rect 25870 5879 25926 5888
rect 26148 5908 26200 5914
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25056 5574 25084 5714
rect 25884 5710 25912 5879
rect 26148 5850 26200 5856
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25608 5234 25636 5646
rect 25976 5234 26004 5646
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25424 4554 25452 5102
rect 25608 4758 25636 5170
rect 26620 5166 26648 5306
rect 26792 5296 26844 5302
rect 26792 5238 26844 5244
rect 25872 5160 25924 5166
rect 25870 5128 25872 5137
rect 26608 5160 26660 5166
rect 25924 5128 25926 5137
rect 26608 5102 26660 5108
rect 26804 5098 26832 5238
rect 25870 5063 25926 5072
rect 26792 5092 26844 5098
rect 26792 5034 26844 5040
rect 26148 5024 26200 5030
rect 26148 4966 26200 4972
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 25596 4752 25648 4758
rect 25596 4694 25648 4700
rect 25412 4548 25464 4554
rect 25412 4490 25464 4496
rect 26160 4486 26188 4966
rect 26252 4826 26280 4966
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26712 4622 26740 4966
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 25228 3528 25280 3534
rect 25504 3528 25556 3534
rect 25228 3470 25280 3476
rect 25502 3496 25504 3505
rect 25556 3496 25558 3505
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24188 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 24540 2202
rect 24188 1114 24540 2150
rect 24596 2106 24624 2382
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 24964 1970 24992 2790
rect 25240 2650 25268 3470
rect 25608 3466 25636 3674
rect 25780 3664 25832 3670
rect 25832 3612 26004 3618
rect 25780 3606 26004 3612
rect 25792 3590 26004 3606
rect 25976 3534 26004 3590
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 25502 3431 25558 3440
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25792 3194 25820 3470
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 26068 3126 26096 3674
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25332 2650 25360 2926
rect 26252 2922 26280 3334
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26240 2916 26292 2922
rect 26240 2858 26292 2864
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 24676 1896 24728 1902
rect 24676 1838 24728 1844
rect 24188 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 24540 1114
rect 24188 1040 24540 1062
rect 24044 870 24164 898
rect 24136 800 24164 870
rect 24688 800 24716 1838
rect 25240 800 25268 2382
rect 25884 1970 25912 2518
rect 25976 2514 26004 2790
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 25872 1964 25924 1970
rect 25872 1906 25924 1912
rect 26068 1562 26096 2382
rect 26160 1970 26188 2382
rect 26148 1964 26200 1970
rect 26148 1906 26200 1912
rect 26056 1556 26108 1562
rect 26056 1498 26108 1504
rect 26332 1352 26384 1358
rect 26332 1294 26384 1300
rect 25780 1284 25832 1290
rect 25780 1226 25832 1232
rect 25792 800 25820 1226
rect 26344 800 26372 1294
rect 26528 1222 26556 2790
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 26700 2304 26752 2310
rect 26700 2246 26752 2252
rect 26712 1970 26740 2246
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 26516 1216 26568 1222
rect 26516 1158 26568 1164
rect 26896 800 26924 2382
rect 26988 1766 27016 2994
rect 27080 2990 27108 6190
rect 27540 5166 27568 6598
rect 29274 6559 29330 6568
rect 28908 6520 28960 6526
rect 28908 6462 28960 6468
rect 28446 5400 28502 5409
rect 28446 5335 28502 5344
rect 28460 5234 28488 5335
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27724 4758 27752 5170
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 28184 5114 28212 5170
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27632 4146 27660 4218
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27632 3942 27660 4082
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27172 3058 27200 3334
rect 27724 3194 27752 3402
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27540 2650 27568 2926
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27816 2514 27844 4966
rect 27908 4758 27936 4966
rect 27896 4752 27948 4758
rect 27896 4694 27948 4700
rect 28000 4078 28028 5102
rect 28184 5086 28856 5114
rect 28828 5030 28856 5086
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 27908 3482 27936 3538
rect 28184 3505 28212 3538
rect 28170 3496 28226 3505
rect 27908 3454 28028 3482
rect 28000 3398 28028 3454
rect 28170 3431 28226 3440
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 27804 2508 27856 2514
rect 27804 2450 27856 2456
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 26976 1760 27028 1766
rect 26976 1702 27028 1708
rect 27448 800 27476 2382
rect 27804 1352 27856 1358
rect 27804 1294 27856 1300
rect 27816 950 27844 1294
rect 27908 1222 27936 3334
rect 28552 3058 28580 4966
rect 28736 3534 28764 4966
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28920 2990 28948 6462
rect 29288 5098 29316 6559
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 29276 5092 29328 5098
rect 29276 5034 29328 5040
rect 29012 5001 29040 5034
rect 29092 5024 29144 5030
rect 28998 4992 29054 5001
rect 29092 4966 29144 4972
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 28998 4927 29054 4936
rect 29104 4622 29132 4966
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28172 2848 28224 2854
rect 28092 2796 28172 2802
rect 28092 2790 28224 2796
rect 28092 2774 28212 2790
rect 27988 1420 28040 1426
rect 27988 1362 28040 1368
rect 27896 1216 27948 1222
rect 27896 1158 27948 1164
rect 27804 944 27856 950
rect 27804 886 27856 892
rect 28000 800 28028 1362
rect 28092 1358 28120 2774
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 28460 1902 28488 2450
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28540 2304 28592 2310
rect 28540 2246 28592 2252
rect 28552 2038 28580 2246
rect 28540 2032 28592 2038
rect 28540 1974 28592 1980
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 28644 1562 28672 2382
rect 28632 1556 28684 1562
rect 28632 1498 28684 1504
rect 29012 1358 29040 4558
rect 29380 3126 29408 4966
rect 29368 3120 29420 3126
rect 29368 3062 29420 3068
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29104 2650 29132 2994
rect 29472 2922 29500 4966
rect 29564 3194 29592 5850
rect 29656 5234 29684 6695
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 30300 5166 30328 6831
rect 31836 6010 32188 7944
rect 34058 7576 34114 7585
rect 34058 7511 34114 7520
rect 32956 6384 33008 6390
rect 32956 6326 33008 6332
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 31836 5958 31858 6010
rect 31910 5958 31922 6010
rect 31974 5958 31986 6010
rect 32038 5958 32050 6010
rect 32102 5958 32114 6010
rect 32166 5958 32188 6010
rect 31576 5568 31628 5574
rect 31576 5510 31628 5516
rect 31208 5296 31260 5302
rect 30838 5264 30894 5273
rect 31208 5238 31260 5244
rect 30838 5199 30840 5208
rect 30892 5199 30894 5208
rect 30840 5170 30892 5176
rect 30288 5160 30340 5166
rect 30380 5160 30432 5166
rect 30288 5102 30340 5108
rect 30378 5128 30380 5137
rect 30432 5128 30434 5137
rect 29644 5092 29696 5098
rect 30378 5063 30434 5072
rect 29644 5034 29696 5040
rect 29656 5001 29684 5034
rect 30472 5024 30524 5030
rect 29642 4992 29698 5001
rect 30472 4966 30524 4972
rect 29642 4927 29698 4936
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29656 3058 29684 4422
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29748 3738 29776 4014
rect 29736 3732 29788 3738
rect 29736 3674 29788 3680
rect 30024 3058 30052 4762
rect 30104 4548 30156 4554
rect 30104 4490 30156 4496
rect 30116 4214 30144 4490
rect 30104 4208 30156 4214
rect 30104 4150 30156 4156
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 29460 2916 29512 2922
rect 29460 2858 29512 2864
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 29092 2304 29144 2310
rect 29092 2246 29144 2252
rect 29104 1970 29132 2246
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 29000 1352 29052 1358
rect 29196 1306 29224 2382
rect 29564 1970 29592 2994
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29920 1964 29972 1970
rect 29920 1906 29972 1912
rect 29000 1294 29052 1300
rect 29104 1278 29224 1306
rect 28540 944 28592 950
rect 28540 886 28592 892
rect 28552 800 28580 886
rect 29104 800 29132 1278
rect 29656 870 29776 898
rect 29656 800 29684 870
rect 3146 0 3202 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 29748 762 29776 870
rect 29932 762 29960 1906
rect 30208 800 30236 2926
rect 30484 2582 30512 4966
rect 31220 3534 31248 5238
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31404 4690 31432 5170
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31312 4049 31340 4082
rect 31298 4040 31354 4049
rect 31298 3975 31354 3984
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31298 3496 31354 3505
rect 31298 3431 31354 3440
rect 31312 3398 31340 3431
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30944 2514 30972 2790
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30300 1902 30328 2246
rect 30288 1896 30340 1902
rect 30288 1838 30340 1844
rect 31036 1562 31064 2382
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31312 1970 31340 2246
rect 31300 1964 31352 1970
rect 31300 1906 31352 1912
rect 31024 1556 31076 1562
rect 31024 1498 31076 1504
rect 31116 1488 31168 1494
rect 31300 1488 31352 1494
rect 31168 1436 31300 1442
rect 31116 1430 31352 1436
rect 31128 1414 31340 1430
rect 30380 1352 30432 1358
rect 30380 1294 30432 1300
rect 29748 734 29960 762
rect 30194 0 30250 800
rect 30392 762 30420 1294
rect 31300 1284 31352 1290
rect 31300 1226 31352 1232
rect 30668 870 30788 898
rect 30668 762 30696 870
rect 30760 800 30788 870
rect 31312 800 31340 1226
rect 31404 1018 31432 3334
rect 31496 3058 31524 4082
rect 31588 3534 31616 5510
rect 31836 4922 32188 5958
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 31836 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 32188 4922
rect 31836 3834 32188 4870
rect 31836 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 32188 3834
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31680 2582 31708 2994
rect 31836 2746 32188 3782
rect 32232 3534 32260 5714
rect 32312 4820 32364 4826
rect 32312 4762 32364 4768
rect 32324 3738 32352 4762
rect 32588 4548 32640 4554
rect 32588 4490 32640 4496
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32218 3088 32274 3097
rect 32218 3023 32274 3032
rect 32312 3052 32364 3058
rect 32232 2990 32260 3023
rect 32312 2994 32364 3000
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 31836 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 32188 2746
rect 31668 2576 31720 2582
rect 31668 2518 31720 2524
rect 31836 2236 32188 2694
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 31836 2180 31864 2236
rect 31920 2180 31944 2236
rect 32000 2180 32024 2236
rect 32080 2180 32104 2236
rect 32160 2180 32188 2236
rect 31836 2156 32188 2180
rect 31836 2100 31864 2156
rect 31920 2100 31944 2156
rect 32000 2100 32024 2156
rect 32080 2100 32104 2156
rect 32160 2100 32188 2156
rect 31836 2076 32188 2100
rect 31836 2020 31864 2076
rect 31920 2020 31944 2076
rect 32000 2020 32024 2076
rect 32080 2020 32104 2076
rect 32160 2020 32188 2076
rect 31836 1996 32188 2020
rect 31836 1940 31864 1996
rect 31920 1940 31944 1996
rect 32000 1940 32024 1996
rect 32080 1940 32104 1996
rect 32160 1940 32188 1996
rect 31836 1658 32188 1940
rect 31836 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 32188 1658
rect 31836 1040 32188 1606
rect 31392 1012 31444 1018
rect 31392 954 31444 960
rect 31864 870 31984 898
rect 31864 800 31892 870
rect 30392 734 30696 762
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 31956 762 31984 870
rect 32232 762 32260 2382
rect 32324 2106 32352 2994
rect 32600 2854 32628 4490
rect 32680 3664 32732 3670
rect 32680 3606 32732 3612
rect 32770 3632 32826 3641
rect 32588 2848 32640 2854
rect 32588 2790 32640 2796
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 2106 32536 2382
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 32496 2100 32548 2106
rect 32496 2042 32548 2048
rect 32404 1896 32456 1902
rect 32404 1838 32456 1844
rect 32416 800 32444 1838
rect 32692 1562 32720 3606
rect 32770 3567 32772 3576
rect 32824 3567 32826 3576
rect 32772 3538 32824 3544
rect 32876 3534 32904 6258
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 32968 2854 32996 6326
rect 33876 5772 33928 5778
rect 33876 5714 33928 5720
rect 33324 5568 33376 5574
rect 33324 5510 33376 5516
rect 33232 3732 33284 3738
rect 33232 3674 33284 3680
rect 33244 3505 33272 3674
rect 33230 3496 33286 3505
rect 33230 3431 33286 3440
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33140 3052 33192 3058
rect 33140 2994 33192 3000
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 33152 2582 33180 2994
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 33048 2304 33100 2310
rect 33048 2246 33100 2252
rect 32680 1556 32732 1562
rect 32680 1498 32732 1504
rect 33060 1426 33088 2246
rect 33048 1420 33100 1426
rect 33048 1362 33100 1368
rect 33244 1358 33272 3130
rect 33336 3058 33364 5510
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 33888 2854 33916 5714
rect 34072 4690 34100 7511
rect 34188 5466 34540 7944
rect 41050 7712 41106 7721
rect 41050 7647 41106 7656
rect 34888 6112 34940 6118
rect 34888 6054 34940 6060
rect 34188 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34540 5466
rect 34060 4684 34112 4690
rect 34060 4626 34112 4632
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 34188 4588 34540 5414
rect 33980 3942 34008 4558
rect 34188 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34540 4588
rect 34188 4508 34540 4532
rect 34188 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34540 4508
rect 34188 4428 34540 4452
rect 34188 4378 34216 4428
rect 34272 4378 34296 4428
rect 34352 4378 34376 4428
rect 34432 4378 34456 4428
rect 34512 4378 34540 4428
rect 34704 4480 34756 4486
rect 34704 4422 34756 4428
rect 34188 4326 34210 4378
rect 34272 4372 34274 4378
rect 34454 4372 34456 4378
rect 34262 4348 34274 4372
rect 34326 4348 34338 4372
rect 34390 4348 34402 4372
rect 34454 4348 34466 4372
rect 34272 4326 34274 4348
rect 34454 4326 34456 4348
rect 34518 4326 34540 4378
rect 34188 4292 34216 4326
rect 34272 4292 34296 4326
rect 34352 4292 34376 4326
rect 34432 4292 34456 4326
rect 34512 4292 34540 4326
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 34188 3290 34540 4292
rect 34716 4146 34744 4422
rect 34796 4276 34848 4282
rect 34796 4218 34848 4224
rect 34808 4146 34836 4218
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34704 4140 34756 4146
rect 34704 4082 34756 4088
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 34624 3890 34652 4082
rect 34808 3942 34836 4082
rect 34796 3936 34848 3942
rect 34624 3862 34744 3890
rect 34796 3878 34848 3884
rect 34188 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34540 3290
rect 34060 3052 34112 3058
rect 34060 2994 34112 3000
rect 33876 2848 33928 2854
rect 33876 2790 33928 2796
rect 34072 2582 34100 2994
rect 34060 2576 34112 2582
rect 34060 2518 34112 2524
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33232 1352 33284 1358
rect 33232 1294 33284 1300
rect 33508 1352 33560 1358
rect 33508 1294 33560 1300
rect 33140 1284 33192 1290
rect 32968 1244 33140 1272
rect 32968 800 32996 1244
rect 33140 1226 33192 1232
rect 33520 800 33548 1294
rect 33612 1222 33640 2382
rect 34188 2202 34540 3238
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 34188 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34540 2202
rect 34060 1964 34112 1970
rect 34060 1906 34112 1912
rect 33600 1216 33652 1222
rect 33600 1158 33652 1164
rect 34072 800 34100 1906
rect 34188 1114 34540 2150
rect 34624 2106 34652 2994
rect 34716 2854 34744 3862
rect 34900 3058 34928 6054
rect 40406 5808 40462 5817
rect 40406 5743 40462 5752
rect 40420 5710 40448 5743
rect 40408 5704 40460 5710
rect 37002 5672 37058 5681
rect 40408 5646 40460 5652
rect 37002 5607 37004 5616
rect 37056 5607 37058 5616
rect 37004 5578 37056 5584
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35072 4752 35124 4758
rect 35072 4694 35124 4700
rect 34980 4140 35032 4146
rect 34980 4082 35032 4088
rect 34992 3194 35020 4082
rect 34980 3188 35032 3194
rect 34980 3130 35032 3136
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34612 2100 34664 2106
rect 34612 2042 34664 2048
rect 34808 1970 34836 2926
rect 35084 2310 35112 4694
rect 35808 3936 35860 3942
rect 35808 3878 35860 3884
rect 35820 2990 35848 3878
rect 35808 2984 35860 2990
rect 35808 2926 35860 2932
rect 35820 2854 35848 2926
rect 35808 2848 35860 2854
rect 35808 2790 35860 2796
rect 35440 2508 35492 2514
rect 35440 2450 35492 2456
rect 35072 2304 35124 2310
rect 35072 2246 35124 2252
rect 34796 1964 34848 1970
rect 34796 1906 34848 1912
rect 34612 1896 34664 1902
rect 34612 1838 34664 1844
rect 34188 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34540 1114
rect 34188 1040 34540 1062
rect 34624 800 34652 1838
rect 35176 870 35296 898
rect 35176 800 35204 870
rect 31956 734 32260 762
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35268 762 35296 870
rect 35452 762 35480 2450
rect 35912 1834 35940 5510
rect 41064 5166 41092 7647
rect 41836 6010 42188 7944
rect 43536 7744 43588 7750
rect 43536 7686 43588 7692
rect 42616 6724 42668 6730
rect 42616 6666 42668 6672
rect 41836 5958 41858 6010
rect 41910 5958 41922 6010
rect 41974 5958 41986 6010
rect 42038 5958 42050 6010
rect 42102 5958 42114 6010
rect 42166 5958 42188 6010
rect 41604 5704 41656 5710
rect 41604 5646 41656 5652
rect 41694 5672 41750 5681
rect 40408 5160 40460 5166
rect 40408 5102 40460 5108
rect 41052 5160 41104 5166
rect 41052 5102 41104 5108
rect 41512 5160 41564 5166
rect 41512 5102 41564 5108
rect 36820 4684 36872 4690
rect 36820 4626 36872 4632
rect 36544 4548 36596 4554
rect 36544 4490 36596 4496
rect 36556 4282 36584 4490
rect 36544 4276 36596 4282
rect 36544 4218 36596 4224
rect 36176 3664 36228 3670
rect 36082 3632 36138 3641
rect 36176 3606 36228 3612
rect 36082 3567 36084 3576
rect 36136 3567 36138 3576
rect 36084 3538 36136 3544
rect 36188 3058 36216 3606
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36636 3052 36688 3058
rect 36636 2994 36688 3000
rect 36648 2106 36676 2994
rect 36740 2938 36768 3130
rect 36832 3058 36860 4626
rect 40420 4010 40448 5102
rect 41524 4826 41552 5102
rect 41512 4820 41564 4826
rect 41512 4762 41564 4768
rect 41236 4616 41288 4622
rect 41236 4558 41288 4564
rect 40408 4004 40460 4010
rect 40408 3946 40460 3952
rect 37004 3936 37056 3942
rect 37004 3878 37056 3884
rect 37016 3194 37044 3878
rect 41248 3738 41276 4558
rect 41236 3732 41288 3738
rect 41236 3674 41288 3680
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 37108 3126 37136 3470
rect 39764 3392 39816 3398
rect 39764 3334 39816 3340
rect 37096 3120 37148 3126
rect 37096 3062 37148 3068
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 37096 2984 37148 2990
rect 36740 2932 37096 2938
rect 36740 2926 37148 2932
rect 36740 2910 37136 2926
rect 39396 2576 39448 2582
rect 39396 2518 39448 2524
rect 39120 2372 39172 2378
rect 39120 2314 39172 2320
rect 39132 2106 39160 2314
rect 39408 2310 39436 2518
rect 39396 2304 39448 2310
rect 39396 2246 39448 2252
rect 39580 2304 39632 2310
rect 39580 2246 39632 2252
rect 36636 2100 36688 2106
rect 36636 2042 36688 2048
rect 39120 2100 39172 2106
rect 39120 2042 39172 2048
rect 39028 1964 39080 1970
rect 39028 1906 39080 1912
rect 36176 1896 36228 1902
rect 36176 1838 36228 1844
rect 37556 1896 37608 1902
rect 37556 1838 37608 1844
rect 35900 1828 35952 1834
rect 35900 1770 35952 1776
rect 35624 1352 35676 1358
rect 35624 1294 35676 1300
rect 35636 1018 35664 1294
rect 36188 1290 36216 1838
rect 37568 1562 37596 1838
rect 37464 1556 37516 1562
rect 37464 1498 37516 1504
rect 37556 1556 37608 1562
rect 37556 1498 37608 1504
rect 37476 1358 37504 1498
rect 37924 1420 37976 1426
rect 37924 1362 37976 1368
rect 37372 1352 37424 1358
rect 37372 1294 37424 1300
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 36176 1284 36228 1290
rect 36176 1226 36228 1232
rect 36268 1284 36320 1290
rect 36268 1226 36320 1232
rect 35716 1216 35768 1222
rect 35716 1158 35768 1164
rect 35624 1012 35676 1018
rect 35624 954 35676 960
rect 35728 800 35756 1158
rect 36280 800 36308 1226
rect 37384 800 37412 1294
rect 37936 800 37964 1362
rect 39040 800 39068 1906
rect 39592 1766 39620 2246
rect 39580 1760 39632 1766
rect 39580 1702 39632 1708
rect 39776 1358 39804 3334
rect 41144 1896 41196 1902
rect 41144 1838 41196 1844
rect 41156 1562 41184 1838
rect 41144 1556 41196 1562
rect 41144 1498 41196 1504
rect 41616 1494 41644 5646
rect 41694 5607 41750 5616
rect 41708 5574 41736 5607
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41836 4922 42188 5958
rect 41836 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 42188 4922
rect 41696 4616 41748 4622
rect 41696 4558 41748 4564
rect 41708 4078 41736 4558
rect 41696 4072 41748 4078
rect 41696 4014 41748 4020
rect 41836 3834 42188 4870
rect 42628 4826 42656 6666
rect 43548 5710 43576 7686
rect 43536 5704 43588 5710
rect 43536 5646 43588 5652
rect 43628 5704 43680 5710
rect 43628 5646 43680 5652
rect 42984 5228 43036 5234
rect 42984 5170 43036 5176
rect 42616 4820 42668 4826
rect 42616 4762 42668 4768
rect 42996 4758 43024 5170
rect 42984 4752 43036 4758
rect 42984 4694 43036 4700
rect 43352 4616 43404 4622
rect 43352 4558 43404 4564
rect 42984 4140 43036 4146
rect 42984 4082 43036 4088
rect 41836 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 42188 3834
rect 41836 2746 42188 3782
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 41836 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 42188 2746
rect 41696 2440 41748 2446
rect 41696 2382 41748 2388
rect 41708 2106 41736 2382
rect 41836 2236 42188 2694
rect 41836 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 42188 2236
rect 41836 2156 42188 2180
rect 41696 2100 41748 2106
rect 41696 2042 41748 2048
rect 41836 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 42188 2156
rect 41836 2076 42188 2100
rect 41836 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 42188 2076
rect 41836 1996 42188 2020
rect 41836 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 42188 1996
rect 41836 1658 42188 1940
rect 42260 1766 42288 3470
rect 42432 3120 42484 3126
rect 42432 3062 42484 3068
rect 42340 2440 42392 2446
rect 42340 2382 42392 2388
rect 42248 1760 42300 1766
rect 42248 1702 42300 1708
rect 41836 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 42188 1658
rect 41604 1488 41656 1494
rect 41604 1430 41656 1436
rect 41236 1420 41288 1426
rect 41236 1362 41288 1368
rect 39764 1352 39816 1358
rect 39764 1294 39816 1300
rect 40776 1352 40828 1358
rect 40776 1294 40828 1300
rect 39580 1284 39632 1290
rect 39580 1226 39632 1232
rect 39592 800 39620 1226
rect 40788 898 40816 1294
rect 40696 870 40816 898
rect 40696 800 40724 870
rect 41248 800 41276 1362
rect 41836 1040 42188 1606
rect 42352 800 42380 2382
rect 42444 1358 42472 3062
rect 42996 1970 43024 4082
rect 43364 2582 43392 4558
rect 43352 2576 43404 2582
rect 43352 2518 43404 2524
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 43076 2372 43128 2378
rect 43076 2314 43128 2320
rect 42892 1964 42944 1970
rect 42892 1906 42944 1912
rect 42984 1964 43036 1970
rect 42984 1906 43036 1912
rect 42904 1358 42932 1906
rect 42984 1828 43036 1834
rect 42984 1770 43036 1776
rect 42432 1352 42484 1358
rect 42432 1294 42484 1300
rect 42892 1352 42944 1358
rect 42892 1294 42944 1300
rect 42996 1000 43024 1770
rect 43088 1426 43116 2314
rect 43076 1420 43128 1426
rect 43076 1362 43128 1368
rect 42904 972 43024 1000
rect 42904 800 42932 972
rect 43456 800 43484 2382
rect 43640 882 43668 5646
rect 44188 5466 44540 7944
rect 48044 7676 48096 7682
rect 48044 7618 48096 7624
rect 46112 6860 46164 6866
rect 46112 6802 46164 6808
rect 45652 6248 45704 6254
rect 45652 6190 45704 6196
rect 44916 6180 44968 6186
rect 44916 6122 44968 6128
rect 44638 5944 44694 5953
rect 44638 5879 44694 5888
rect 44652 5710 44680 5879
rect 44928 5778 44956 6122
rect 45560 6112 45612 6118
rect 45560 6054 45612 6060
rect 44916 5772 44968 5778
rect 44916 5714 44968 5720
rect 45572 5710 45600 6054
rect 45664 5710 45692 6190
rect 44640 5704 44692 5710
rect 44640 5646 44692 5652
rect 45560 5704 45612 5710
rect 45560 5646 45612 5652
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 45928 5568 45980 5574
rect 45928 5510 45980 5516
rect 46018 5536 46074 5545
rect 44188 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 44540 5466
rect 44088 5160 44140 5166
rect 44086 5128 44088 5137
rect 44140 5128 44142 5137
rect 44086 5063 44142 5072
rect 44188 4588 44540 5414
rect 45940 5234 45968 5510
rect 46018 5471 46074 5480
rect 45928 5228 45980 5234
rect 45928 5170 45980 5176
rect 46032 5166 46060 5471
rect 44640 5160 44692 5166
rect 44640 5102 44692 5108
rect 45376 5160 45428 5166
rect 45376 5102 45428 5108
rect 46020 5160 46072 5166
rect 46020 5102 46072 5108
rect 44188 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 44540 4588
rect 44188 4508 44540 4532
rect 43904 4480 43956 4486
rect 43904 4422 43956 4428
rect 44188 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 44540 4508
rect 44188 4428 44540 4452
rect 43916 4146 43944 4422
rect 44188 4378 44216 4428
rect 44272 4378 44296 4428
rect 44352 4378 44376 4428
rect 44432 4378 44456 4428
rect 44512 4378 44540 4428
rect 44188 4326 44210 4378
rect 44272 4372 44274 4378
rect 44454 4372 44456 4378
rect 44262 4348 44274 4372
rect 44326 4348 44338 4372
rect 44390 4348 44402 4372
rect 44454 4348 44466 4372
rect 44272 4326 44274 4348
rect 44454 4326 44456 4348
rect 44518 4326 44540 4378
rect 44188 4292 44216 4326
rect 44272 4292 44296 4326
rect 44352 4292 44376 4326
rect 44432 4292 44456 4326
rect 44512 4292 44540 4326
rect 43904 4140 43956 4146
rect 43904 4082 43956 4088
rect 44188 3290 44540 4292
rect 44652 3602 44680 5102
rect 45008 5024 45060 5030
rect 44730 4992 44786 5001
rect 45008 4966 45060 4972
rect 45100 5024 45152 5030
rect 45100 4966 45152 4972
rect 44730 4927 44786 4936
rect 44744 4758 44772 4927
rect 45020 4758 45048 4966
rect 45112 4826 45140 4966
rect 45100 4820 45152 4826
rect 45100 4762 45152 4768
rect 44732 4752 44784 4758
rect 44732 4694 44784 4700
rect 45008 4752 45060 4758
rect 45008 4694 45060 4700
rect 44640 3596 44692 3602
rect 44640 3538 44692 3544
rect 45388 3466 45416 5102
rect 46124 5030 46152 6802
rect 46388 6520 46440 6526
rect 46388 6462 46440 6468
rect 46400 5710 46428 6462
rect 47032 6180 47084 6186
rect 47032 6122 47084 6128
rect 47044 5710 47072 6122
rect 47492 5908 47544 5914
rect 47492 5850 47544 5856
rect 47504 5710 47532 5850
rect 46388 5704 46440 5710
rect 46388 5646 46440 5652
rect 47032 5704 47084 5710
rect 47032 5646 47084 5652
rect 47492 5704 47544 5710
rect 47492 5646 47544 5652
rect 47400 5568 47452 5574
rect 47400 5510 47452 5516
rect 46216 5358 46520 5386
rect 46216 5302 46244 5358
rect 46492 5302 46520 5358
rect 46204 5296 46256 5302
rect 46204 5238 46256 5244
rect 46480 5296 46532 5302
rect 46480 5238 46532 5244
rect 46296 5228 46348 5234
rect 46296 5170 46348 5176
rect 46112 5024 46164 5030
rect 46112 4966 46164 4972
rect 46308 4622 46336 5170
rect 46388 5160 46440 5166
rect 46388 5102 46440 5108
rect 46296 4616 46348 4622
rect 46296 4558 46348 4564
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 45376 3460 45428 3466
rect 45376 3402 45428 3408
rect 44916 3392 44968 3398
rect 44916 3334 44968 3340
rect 44188 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 44540 3290
rect 44188 2202 44540 3238
rect 44824 2916 44876 2922
rect 44824 2858 44876 2864
rect 44732 2576 44784 2582
rect 44732 2518 44784 2524
rect 44188 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 44540 2202
rect 43996 1284 44048 1290
rect 43996 1226 44048 1232
rect 43628 876 43680 882
rect 43628 818 43680 824
rect 44008 800 44036 1226
rect 44188 1114 44540 2150
rect 44744 1358 44772 2518
rect 44836 1748 44864 2858
rect 44928 2854 44956 3334
rect 45940 3058 45968 4422
rect 45928 3052 45980 3058
rect 45928 2994 45980 3000
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44928 1902 44956 2790
rect 45560 2440 45612 2446
rect 45560 2382 45612 2388
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 45376 1964 45428 1970
rect 45376 1906 45428 1912
rect 44916 1896 44968 1902
rect 44916 1838 44968 1844
rect 44836 1720 44956 1748
rect 44824 1420 44876 1426
rect 44824 1362 44876 1368
rect 44732 1352 44784 1358
rect 44732 1294 44784 1300
rect 44188 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 44540 1114
rect 44188 1040 44540 1062
rect 44560 870 44680 898
rect 44560 800 44588 870
rect 35268 734 35480 762
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 44652 762 44680 870
rect 44836 762 44864 1362
rect 44928 1358 44956 1720
rect 45388 1562 45416 1906
rect 45572 1562 45600 2382
rect 45652 1964 45704 1970
rect 45652 1906 45704 1912
rect 45376 1556 45428 1562
rect 45376 1498 45428 1504
rect 45560 1556 45612 1562
rect 45560 1498 45612 1504
rect 44916 1352 44968 1358
rect 44916 1294 44968 1300
rect 45100 1284 45152 1290
rect 45100 1226 45152 1232
rect 45112 800 45140 1226
rect 45664 800 45692 1906
rect 46216 1902 46244 2382
rect 46400 2378 46428 5102
rect 47044 5098 47256 5114
rect 47032 5092 47256 5098
rect 47084 5086 47256 5092
rect 47228 5080 47256 5086
rect 47308 5092 47360 5098
rect 47228 5052 47308 5080
rect 47032 5034 47084 5040
rect 47308 5034 47360 5040
rect 47412 5030 47440 5510
rect 48056 5166 48084 7618
rect 48872 6792 48924 6798
rect 48872 6734 48924 6740
rect 48228 6384 48280 6390
rect 48228 6326 48280 6332
rect 48136 6248 48188 6254
rect 48136 6190 48188 6196
rect 48148 5914 48176 6190
rect 48136 5908 48188 5914
rect 48136 5850 48188 5856
rect 48240 5710 48268 6326
rect 48884 5914 48912 6734
rect 51724 6520 51776 6526
rect 51724 6462 51776 6468
rect 51080 6316 51132 6322
rect 51080 6258 51132 6264
rect 51092 6186 51120 6258
rect 51080 6180 51132 6186
rect 51080 6122 51132 6128
rect 49514 6080 49570 6089
rect 49514 6015 49570 6024
rect 48872 5908 48924 5914
rect 48872 5850 48924 5856
rect 48228 5704 48280 5710
rect 48228 5646 48280 5652
rect 49528 5642 49556 6015
rect 51736 5778 51764 6462
rect 51836 6010 52188 7944
rect 52276 7812 52328 7818
rect 52276 7754 52328 7760
rect 51836 5958 51858 6010
rect 51910 5958 51922 6010
rect 51974 5958 51986 6010
rect 52038 5958 52050 6010
rect 52102 5958 52114 6010
rect 52166 5958 52188 6010
rect 49792 5772 49844 5778
rect 49792 5714 49844 5720
rect 51724 5772 51776 5778
rect 51724 5714 51776 5720
rect 49516 5636 49568 5642
rect 49516 5578 49568 5584
rect 49804 5166 49832 5714
rect 50436 5704 50488 5710
rect 50436 5646 50488 5652
rect 51264 5704 51316 5710
rect 51264 5646 51316 5652
rect 47492 5160 47544 5166
rect 48044 5160 48096 5166
rect 47492 5102 47544 5108
rect 47582 5128 47638 5137
rect 47124 5024 47176 5030
rect 47124 4966 47176 4972
rect 47400 5024 47452 5030
rect 47400 4966 47452 4972
rect 46662 4856 46718 4865
rect 46662 4791 46718 4800
rect 46676 4622 46704 4791
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 46664 4616 46716 4622
rect 46664 4558 46716 4564
rect 46572 4548 46624 4554
rect 46572 4490 46624 4496
rect 46584 4434 46612 4490
rect 46756 4480 46808 4486
rect 46584 4428 46756 4434
rect 46584 4422 46808 4428
rect 46584 4406 46796 4422
rect 47044 4146 47072 4626
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 47032 4004 47084 4010
rect 47032 3946 47084 3952
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 46860 1970 46888 2246
rect 47044 2106 47072 3946
rect 47136 3058 47164 4966
rect 47504 4282 47532 5102
rect 48044 5102 48096 5108
rect 49148 5160 49200 5166
rect 49148 5102 49200 5108
rect 49792 5160 49844 5166
rect 49792 5102 49844 5108
rect 47582 5063 47638 5072
rect 47596 4282 47624 5063
rect 48964 4548 49016 4554
rect 48964 4490 49016 4496
rect 47492 4276 47544 4282
rect 47492 4218 47544 4224
rect 47584 4276 47636 4282
rect 47584 4218 47636 4224
rect 48976 4146 49004 4490
rect 49056 4480 49108 4486
rect 49056 4422 49108 4428
rect 48964 4140 49016 4146
rect 48964 4082 49016 4088
rect 47400 3936 47452 3942
rect 47400 3878 47452 3884
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 47308 2440 47360 2446
rect 47308 2382 47360 2388
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47032 2100 47084 2106
rect 47032 2042 47084 2048
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46020 1896 46072 1902
rect 46020 1838 46072 1844
rect 46204 1896 46256 1902
rect 46204 1838 46256 1844
rect 46032 1222 46060 1838
rect 47228 1562 47256 2314
rect 47216 1556 47268 1562
rect 47216 1498 47268 1504
rect 46204 1420 46256 1426
rect 46204 1362 46256 1368
rect 46020 1216 46072 1222
rect 46020 1158 46072 1164
rect 46216 800 46244 1362
rect 47320 800 47348 2382
rect 47412 1358 47440 3878
rect 47858 3360 47914 3369
rect 47858 3295 47914 3304
rect 47584 2848 47636 2854
rect 47584 2790 47636 2796
rect 47596 1970 47624 2790
rect 47872 2514 47900 3295
rect 49068 3058 49096 4422
rect 49160 3670 49188 5102
rect 49332 5024 49384 5030
rect 49332 4966 49384 4972
rect 49344 4758 49372 4966
rect 49332 4752 49384 4758
rect 49332 4694 49384 4700
rect 49148 3664 49200 3670
rect 49148 3606 49200 3612
rect 49056 3052 49108 3058
rect 49056 2994 49108 3000
rect 50068 2916 50120 2922
rect 50068 2858 50120 2864
rect 47860 2508 47912 2514
rect 47860 2450 47912 2456
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 48056 2106 48084 2450
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 48044 2100 48096 2106
rect 48044 2042 48096 2048
rect 47584 1964 47636 1970
rect 47584 1906 47636 1912
rect 47860 1896 47912 1902
rect 47860 1838 47912 1844
rect 47400 1352 47452 1358
rect 47400 1294 47452 1300
rect 47872 800 47900 1838
rect 49068 1272 49096 2382
rect 49424 2304 49476 2310
rect 49424 2246 49476 2252
rect 49516 2304 49568 2310
rect 49516 2246 49568 2252
rect 49436 1358 49464 2246
rect 49528 1970 49556 2246
rect 49516 1964 49568 1970
rect 49516 1906 49568 1912
rect 49608 1420 49660 1426
rect 49608 1362 49660 1368
rect 49424 1352 49476 1358
rect 49424 1294 49476 1300
rect 48976 1244 49096 1272
rect 48976 800 49004 1244
rect 49620 898 49648 1362
rect 50080 1358 50108 2858
rect 50448 1834 50476 5646
rect 51276 4010 51304 5646
rect 51836 4922 52188 5958
rect 52288 5710 52316 7754
rect 53288 6248 53340 6254
rect 53288 6190 53340 6196
rect 53300 5914 53328 6190
rect 53288 5908 53340 5914
rect 53288 5850 53340 5856
rect 52276 5704 52328 5710
rect 52920 5704 52972 5710
rect 52276 5646 52328 5652
rect 52748 5664 52920 5692
rect 52368 5636 52420 5642
rect 52368 5578 52420 5584
rect 52380 5234 52408 5578
rect 52552 5568 52604 5574
rect 52552 5510 52604 5516
rect 52368 5228 52420 5234
rect 52368 5170 52420 5176
rect 51836 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 52188 4922
rect 51540 4684 51592 4690
rect 51540 4626 51592 4632
rect 51552 4282 51580 4626
rect 51540 4276 51592 4282
rect 51540 4218 51592 4224
rect 51264 4004 51316 4010
rect 51264 3946 51316 3952
rect 51836 3834 52188 4870
rect 51836 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 52188 3834
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 51184 2582 51212 3470
rect 51836 2746 52188 3782
rect 52564 3602 52592 5510
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52644 2848 52696 2854
rect 52644 2790 52696 2796
rect 51836 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 52188 2746
rect 51172 2576 51224 2582
rect 51172 2518 51224 2524
rect 51836 2236 52188 2694
rect 51836 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 52188 2236
rect 51836 2156 52188 2180
rect 51836 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 52188 2156
rect 51836 2076 52188 2100
rect 51836 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 52188 2076
rect 51836 1996 52188 2020
rect 51836 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 52188 1996
rect 51264 1896 51316 1902
rect 51264 1838 51316 1844
rect 50436 1828 50488 1834
rect 50436 1770 50488 1776
rect 51276 1562 51304 1838
rect 51836 1658 52188 1940
rect 51836 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 52188 1658
rect 51264 1556 51316 1562
rect 51264 1498 51316 1504
rect 50068 1352 50120 1358
rect 50068 1294 50120 1300
rect 50620 1352 50672 1358
rect 50620 1294 50672 1300
rect 49528 870 49648 898
rect 49528 800 49556 870
rect 50632 800 50660 1294
rect 51172 1284 51224 1290
rect 51172 1226 51224 1232
rect 51184 800 51212 1226
rect 51836 1040 52188 1606
rect 52656 1358 52684 2790
rect 52748 1834 52776 5664
rect 52920 5646 52972 5652
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 53012 5636 53064 5642
rect 53012 5578 53064 5584
rect 53024 5234 53052 5578
rect 53116 5234 53420 5250
rect 53012 5228 53064 5234
rect 53012 5170 53064 5176
rect 53104 5228 53420 5234
rect 53156 5222 53420 5228
rect 53104 5170 53156 5176
rect 53392 5166 53420 5222
rect 53288 5160 53340 5166
rect 53288 5102 53340 5108
rect 53380 5160 53432 5166
rect 53380 5102 53432 5108
rect 52920 5024 52972 5030
rect 52920 4966 52972 4972
rect 52932 3058 52960 4966
rect 53300 4282 53328 5102
rect 53288 4276 53340 4282
rect 53288 4218 53340 4224
rect 52920 3052 52972 3058
rect 52920 2994 52972 3000
rect 53104 2848 53156 2854
rect 53104 2790 53156 2796
rect 53116 1970 53144 2790
rect 53852 2530 53880 5646
rect 54188 5466 54540 7944
rect 59196 7800 59224 8024
rect 59572 7857 59600 8024
rect 59188 7772 59224 7800
rect 59558 7848 59614 7857
rect 59558 7783 59614 7792
rect 60740 7812 60792 7818
rect 55588 7676 55640 7682
rect 55588 7618 55640 7624
rect 54852 7608 54904 7614
rect 54680 7556 54852 7562
rect 54680 7550 54904 7556
rect 54680 7534 54892 7550
rect 54680 7478 54708 7534
rect 54668 7472 54720 7478
rect 54668 7414 54720 7420
rect 54668 6928 54720 6934
rect 54668 6870 54720 6876
rect 54680 5574 54708 6870
rect 54852 6384 54904 6390
rect 54852 6326 54904 6332
rect 54864 5574 54892 6326
rect 55220 5772 55272 5778
rect 55220 5714 55272 5720
rect 54668 5568 54720 5574
rect 54668 5510 54720 5516
rect 54852 5568 54904 5574
rect 54852 5510 54904 5516
rect 54188 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 54540 5466
rect 54188 4588 54540 5414
rect 54576 5228 54628 5234
rect 54576 5170 54628 5176
rect 54944 5228 54996 5234
rect 54944 5170 54996 5176
rect 55036 5228 55088 5234
rect 55036 5170 55088 5176
rect 54588 5114 54616 5170
rect 54588 5086 54800 5114
rect 54772 5030 54800 5086
rect 54668 5024 54720 5030
rect 54668 4966 54720 4972
rect 54760 5024 54812 5030
rect 54760 4966 54812 4972
rect 54188 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 54540 4588
rect 54188 4508 54540 4532
rect 54188 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 54540 4508
rect 54188 4428 54540 4452
rect 54188 4378 54216 4428
rect 54272 4378 54296 4428
rect 54352 4378 54376 4428
rect 54432 4378 54456 4428
rect 54512 4378 54540 4428
rect 54188 4326 54210 4378
rect 54272 4372 54274 4378
rect 54454 4372 54456 4378
rect 54262 4348 54274 4372
rect 54326 4348 54338 4372
rect 54390 4348 54402 4372
rect 54454 4348 54466 4372
rect 54272 4326 54274 4348
rect 54454 4326 54456 4348
rect 54518 4326 54540 4378
rect 54188 4292 54216 4326
rect 54272 4292 54296 4326
rect 54352 4292 54376 4326
rect 54432 4292 54456 4326
rect 54512 4292 54540 4326
rect 54188 3290 54540 4292
rect 54188 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 54540 3290
rect 53932 3052 53984 3058
rect 53932 2994 53984 3000
rect 53944 2582 53972 2994
rect 53760 2502 53880 2530
rect 53932 2576 53984 2582
rect 53932 2518 53984 2524
rect 54024 2576 54076 2582
rect 54024 2518 54076 2524
rect 53760 2378 53788 2502
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53932 2440 53984 2446
rect 53932 2382 53984 2388
rect 53748 2372 53800 2378
rect 53748 2314 53800 2320
rect 53104 1964 53156 1970
rect 53104 1906 53156 1912
rect 52920 1896 52972 1902
rect 52840 1856 52920 1884
rect 52736 1828 52788 1834
rect 52736 1770 52788 1776
rect 52644 1352 52696 1358
rect 52644 1294 52696 1300
rect 52276 1216 52328 1222
rect 52276 1158 52328 1164
rect 52288 800 52316 1158
rect 52840 800 52868 1856
rect 52920 1838 52972 1844
rect 53852 1358 53880 2382
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 53944 800 53972 2382
rect 54036 2106 54064 2518
rect 54188 2202 54540 3238
rect 54680 3058 54708 4966
rect 54956 4690 54984 5170
rect 54852 4684 54904 4690
rect 54852 4626 54904 4632
rect 54944 4684 54996 4690
rect 54944 4626 54996 4632
rect 54864 4570 54892 4626
rect 55048 4570 55076 5170
rect 55232 4706 55260 5714
rect 55600 5574 55628 7618
rect 59188 7449 59216 7772
rect 60740 7754 60792 7760
rect 61660 7812 61712 7818
rect 61660 7754 61712 7760
rect 60752 7546 60780 7754
rect 60740 7540 60792 7546
rect 60740 7482 60792 7488
rect 59174 7440 59230 7449
rect 59174 7375 59230 7384
rect 60740 7336 60792 7342
rect 60740 7278 60792 7284
rect 59084 7200 59136 7206
rect 59084 7142 59136 7148
rect 55772 6996 55824 7002
rect 55772 6938 55824 6944
rect 55784 6526 55812 6938
rect 55864 6860 55916 6866
rect 55864 6802 55916 6808
rect 55876 6526 55904 6802
rect 55772 6520 55824 6526
rect 55772 6462 55824 6468
rect 55864 6520 55916 6526
rect 55864 6462 55916 6468
rect 56506 6352 56562 6361
rect 56506 6287 56562 6296
rect 55770 6216 55826 6225
rect 55770 6151 55826 6160
rect 55680 6112 55732 6118
rect 55680 6054 55732 6060
rect 55692 5692 55720 6054
rect 55784 5817 55812 6151
rect 55864 6112 55916 6118
rect 55864 6054 55916 6060
rect 55876 5846 55904 6054
rect 55864 5840 55916 5846
rect 55770 5808 55826 5817
rect 55864 5782 55916 5788
rect 56520 5778 56548 6287
rect 57428 6248 57480 6254
rect 57428 6190 57480 6196
rect 57520 6248 57572 6254
rect 57520 6190 57572 6196
rect 57440 5914 57468 6190
rect 57532 6089 57560 6190
rect 57518 6080 57574 6089
rect 57518 6015 57574 6024
rect 58162 6080 58218 6089
rect 58162 6015 58218 6024
rect 57428 5908 57480 5914
rect 57428 5850 57480 5856
rect 58176 5778 58204 6015
rect 55770 5743 55826 5752
rect 56508 5772 56560 5778
rect 56508 5714 56560 5720
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 58164 5772 58216 5778
rect 58164 5714 58216 5720
rect 56416 5704 56468 5710
rect 55692 5664 56364 5692
rect 56336 5574 56364 5664
rect 56416 5646 56468 5652
rect 55588 5568 55640 5574
rect 56232 5568 56284 5574
rect 55588 5510 55640 5516
rect 55862 5536 55918 5545
rect 56232 5510 56284 5516
rect 56324 5568 56376 5574
rect 56324 5510 56376 5516
rect 55862 5471 55918 5480
rect 55876 5137 55904 5471
rect 55862 5128 55918 5137
rect 55862 5063 55918 5072
rect 54864 4542 55076 4570
rect 55140 4678 55260 4706
rect 55140 4298 55168 4678
rect 55496 4480 55548 4486
rect 55496 4422 55548 4428
rect 55140 4270 55352 4298
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 55220 2848 55272 2854
rect 55220 2790 55272 2796
rect 55036 2372 55088 2378
rect 55036 2314 55088 2320
rect 54760 2304 54812 2310
rect 54760 2246 54812 2252
rect 54188 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 54540 2202
rect 54024 2100 54076 2106
rect 54024 2042 54076 2048
rect 54188 1114 54540 2150
rect 54772 1970 54800 2246
rect 55048 2106 55076 2314
rect 55036 2100 55088 2106
rect 55036 2042 55088 2048
rect 54760 1964 54812 1970
rect 54760 1906 54812 1912
rect 55232 1358 55260 2790
rect 55324 2514 55352 4270
rect 55508 4146 55536 4422
rect 55496 4140 55548 4146
rect 55496 4082 55548 4088
rect 55864 3596 55916 3602
rect 55864 3538 55916 3544
rect 55312 2508 55364 2514
rect 55312 2450 55364 2456
rect 55588 1896 55640 1902
rect 55588 1838 55640 1844
rect 55220 1352 55272 1358
rect 55220 1294 55272 1300
rect 54576 1284 54628 1290
rect 54576 1226 54628 1232
rect 54188 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 54540 1114
rect 54188 1040 54540 1062
rect 54588 898 54616 1226
rect 54496 870 54616 898
rect 54496 800 54524 870
rect 55600 800 55628 1838
rect 55876 1834 55904 3538
rect 56244 3058 56272 5510
rect 56428 5166 56456 5646
rect 56416 5160 56468 5166
rect 56416 5102 56468 5108
rect 57808 3058 57836 5714
rect 59096 5302 59124 7142
rect 60464 7132 60516 7138
rect 60464 7074 60516 7080
rect 59634 7032 59690 7041
rect 59634 6967 59690 6976
rect 59452 5772 59504 5778
rect 59452 5714 59504 5720
rect 59084 5296 59136 5302
rect 59084 5238 59136 5244
rect 59464 3058 59492 5714
rect 59648 5574 59676 6967
rect 60476 6254 60504 7074
rect 60556 6860 60608 6866
rect 60556 6802 60608 6808
rect 60568 6746 60596 6802
rect 60568 6718 60688 6746
rect 60660 6254 60688 6718
rect 60464 6248 60516 6254
rect 60464 6190 60516 6196
rect 60648 6248 60700 6254
rect 60648 6190 60700 6196
rect 60752 5710 60780 7278
rect 61016 6928 61068 6934
rect 60844 6876 61016 6882
rect 60844 6870 61068 6876
rect 60844 6854 61056 6870
rect 61384 6860 61436 6866
rect 60844 6458 60872 6854
rect 61384 6802 61436 6808
rect 61396 6662 61424 6802
rect 61384 6656 61436 6662
rect 61384 6598 61436 6604
rect 60832 6452 60884 6458
rect 60832 6394 60884 6400
rect 61016 6452 61068 6458
rect 61016 6394 61068 6400
rect 61028 6338 61056 6394
rect 60844 6310 61056 6338
rect 60844 5914 60872 6310
rect 60832 5908 60884 5914
rect 60832 5850 60884 5856
rect 61672 5778 61700 7754
rect 61836 6010 62188 7944
rect 62948 7880 63000 7886
rect 62948 7822 63000 7828
rect 62764 7744 62816 7750
rect 62764 7686 62816 7692
rect 62856 7744 62908 7750
rect 62856 7686 62908 7692
rect 62776 7478 62804 7686
rect 62764 7472 62816 7478
rect 62764 7414 62816 7420
rect 62672 7268 62724 7274
rect 62672 7210 62724 7216
rect 61836 5958 61858 6010
rect 61910 5958 61922 6010
rect 61974 5958 61986 6010
rect 62038 5958 62050 6010
rect 62102 5958 62114 6010
rect 62166 5958 62188 6010
rect 61660 5772 61712 5778
rect 61660 5714 61712 5720
rect 60740 5704 60792 5710
rect 60740 5646 60792 5652
rect 60924 5636 60976 5642
rect 60924 5578 60976 5584
rect 61108 5636 61160 5642
rect 61108 5578 61160 5584
rect 59636 5568 59688 5574
rect 60936 5545 60964 5578
rect 59636 5510 59688 5516
rect 60922 5536 60978 5545
rect 60922 5471 60978 5480
rect 61016 5296 61068 5302
rect 61016 5238 61068 5244
rect 61028 4826 61056 5238
rect 61016 4820 61068 4826
rect 61016 4762 61068 4768
rect 61016 4616 61068 4622
rect 61016 4558 61068 4564
rect 60924 4548 60976 4554
rect 60924 4490 60976 4496
rect 60740 4140 60792 4146
rect 60740 4082 60792 4088
rect 56232 3052 56284 3058
rect 56232 2994 56284 3000
rect 57796 3052 57848 3058
rect 57796 2994 57848 3000
rect 59452 3052 59504 3058
rect 59452 2994 59504 3000
rect 56416 2848 56468 2854
rect 56416 2790 56468 2796
rect 57980 2848 58032 2854
rect 57980 2790 58032 2796
rect 60372 2848 60424 2854
rect 60372 2790 60424 2796
rect 56428 1970 56456 2790
rect 57336 2440 57388 2446
rect 57336 2382 57388 2388
rect 56692 2372 56744 2378
rect 56692 2314 56744 2320
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 56140 1896 56192 1902
rect 56140 1838 56192 1844
rect 55864 1828 55916 1834
rect 55864 1770 55916 1776
rect 56152 800 56180 1838
rect 56704 1358 56732 2314
rect 57244 1760 57296 1766
rect 57244 1702 57296 1708
rect 57256 1358 57284 1702
rect 56692 1352 56744 1358
rect 56692 1294 56744 1300
rect 57244 1352 57296 1358
rect 57244 1294 57296 1300
rect 57348 1170 57376 2382
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 57900 1970 57928 2246
rect 57888 1964 57940 1970
rect 57888 1906 57940 1912
rect 57992 1358 58020 2790
rect 59360 1896 59412 1902
rect 59360 1838 59412 1844
rect 59372 1358 59400 1838
rect 59452 1420 59504 1426
rect 59452 1362 59504 1368
rect 57980 1352 58032 1358
rect 57980 1294 58032 1300
rect 59360 1352 59412 1358
rect 59360 1294 59412 1300
rect 57796 1284 57848 1290
rect 57796 1226 57848 1232
rect 58900 1284 58952 1290
rect 58900 1226 58952 1232
rect 57256 1142 57376 1170
rect 57256 800 57284 1142
rect 57808 800 57836 1226
rect 58912 800 58940 1226
rect 59464 800 59492 1362
rect 60384 1358 60412 2790
rect 60752 2378 60780 4082
rect 60936 4010 60964 4490
rect 61028 4185 61056 4558
rect 61120 4486 61148 5578
rect 61200 5568 61252 5574
rect 61200 5510 61252 5516
rect 61108 4480 61160 4486
rect 61108 4422 61160 4428
rect 61014 4176 61070 4185
rect 61014 4111 61070 4120
rect 60924 4004 60976 4010
rect 60924 3946 60976 3952
rect 61212 3058 61240 5510
rect 61292 5228 61344 5234
rect 61292 5170 61344 5176
rect 61304 4706 61332 5170
rect 61836 4922 62188 5958
rect 62580 5908 62632 5914
rect 62580 5850 62632 5856
rect 62592 5778 62620 5850
rect 62580 5772 62632 5778
rect 62580 5714 62632 5720
rect 61836 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 62188 4922
rect 61304 4678 61424 4706
rect 61304 4622 61332 4678
rect 61292 4616 61344 4622
rect 61292 4558 61344 4564
rect 61396 3466 61424 4678
rect 61476 4616 61528 4622
rect 61476 4558 61528 4564
rect 61488 4185 61516 4558
rect 61474 4176 61530 4185
rect 61474 4111 61530 4120
rect 61476 4072 61528 4078
rect 61476 4014 61528 4020
rect 61384 3460 61436 3466
rect 61384 3402 61436 3408
rect 61200 3052 61252 3058
rect 61200 2994 61252 3000
rect 61384 2848 61436 2854
rect 61384 2790 61436 2796
rect 60740 2372 60792 2378
rect 60740 2314 60792 2320
rect 61016 2372 61068 2378
rect 61016 2314 61068 2320
rect 60556 1896 60608 1902
rect 60556 1838 60608 1844
rect 60372 1352 60424 1358
rect 60372 1294 60424 1300
rect 60568 800 60596 1838
rect 61028 1562 61056 2314
rect 61396 1970 61424 2790
rect 61488 2106 61516 4014
rect 61836 3834 62188 4870
rect 62684 4282 62712 7210
rect 62868 6118 62896 7686
rect 62960 6594 62988 7822
rect 63420 7682 63448 10286
rect 63408 7676 63460 7682
rect 63408 7618 63460 7624
rect 63512 7410 63540 11727
rect 63500 7404 63552 7410
rect 63500 7346 63552 7352
rect 63498 7304 63554 7313
rect 63498 7239 63554 7248
rect 62948 6588 63000 6594
rect 62948 6530 63000 6536
rect 63408 6452 63460 6458
rect 63408 6394 63460 6400
rect 63420 6118 63448 6394
rect 62856 6112 62908 6118
rect 62762 6080 62818 6089
rect 63408 6112 63460 6118
rect 62856 6054 62908 6060
rect 63130 6080 63186 6089
rect 62762 6015 62818 6024
rect 63408 6054 63460 6060
rect 63130 6015 63186 6024
rect 62776 5914 62804 6015
rect 62764 5908 62816 5914
rect 62764 5850 62816 5856
rect 62946 5808 63002 5817
rect 62946 5743 63002 5752
rect 62960 5710 62988 5743
rect 62948 5704 63000 5710
rect 62948 5646 63000 5652
rect 63144 5409 63172 6015
rect 63408 5908 63460 5914
rect 63408 5850 63460 5856
rect 63420 5817 63448 5850
rect 63406 5808 63462 5817
rect 63406 5743 63462 5752
rect 63316 5568 63368 5574
rect 63236 5516 63316 5522
rect 63236 5510 63368 5516
rect 63236 5494 63356 5510
rect 63130 5400 63186 5409
rect 63130 5335 63186 5344
rect 62856 5296 62908 5302
rect 62856 5238 62908 5244
rect 62764 4820 62816 4826
rect 62764 4762 62816 4768
rect 62672 4276 62724 4282
rect 62672 4218 62724 4224
rect 62776 4010 62804 4762
rect 62868 4554 62896 5238
rect 62856 4548 62908 4554
rect 62856 4490 62908 4496
rect 62764 4004 62816 4010
rect 62764 3946 62816 3952
rect 61836 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 62188 3834
rect 61836 2746 62188 3782
rect 63236 3058 63264 5494
rect 63406 5400 63462 5409
rect 63406 5335 63462 5344
rect 63420 4865 63448 5335
rect 63512 5030 63540 7239
rect 63604 6361 63632 25774
rect 63684 25764 63736 25770
rect 63684 25706 63736 25712
rect 63696 6798 63724 25706
rect 63788 16561 63816 29582
rect 63774 16552 63830 16561
rect 63774 16487 63830 16496
rect 63776 16448 63828 16454
rect 63776 16390 63828 16396
rect 63788 12050 63816 16390
rect 63880 12170 63908 45222
rect 63868 12164 63920 12170
rect 63868 12106 63920 12112
rect 63788 12022 63908 12050
rect 63776 11892 63828 11898
rect 63776 11834 63828 11840
rect 63684 6792 63736 6798
rect 63684 6734 63736 6740
rect 63684 6452 63736 6458
rect 63684 6394 63736 6400
rect 63590 6352 63646 6361
rect 63590 6287 63646 6296
rect 63592 5636 63644 5642
rect 63592 5578 63644 5584
rect 63604 5370 63632 5578
rect 63592 5364 63644 5370
rect 63592 5306 63644 5312
rect 63500 5024 63552 5030
rect 63500 4966 63552 4972
rect 63406 4856 63462 4865
rect 63406 4791 63462 4800
rect 63590 4856 63646 4865
rect 63590 4791 63646 4800
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 63604 2990 63632 4791
rect 63592 2984 63644 2990
rect 63592 2926 63644 2932
rect 63040 2848 63092 2854
rect 63040 2790 63092 2796
rect 61836 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 62188 2746
rect 61836 2236 62188 2694
rect 62304 2440 62356 2446
rect 62304 2382 62356 2388
rect 61836 2180 61864 2236
rect 61920 2180 61944 2236
rect 62000 2180 62024 2236
rect 62080 2180 62104 2236
rect 62160 2180 62188 2236
rect 61836 2156 62188 2180
rect 61476 2100 61528 2106
rect 61476 2042 61528 2048
rect 61836 2100 61864 2156
rect 61920 2100 61944 2156
rect 62000 2100 62024 2156
rect 62080 2100 62104 2156
rect 62160 2100 62188 2156
rect 61836 2076 62188 2100
rect 61836 2020 61864 2076
rect 61920 2020 61944 2076
rect 62000 2020 62024 2076
rect 62080 2020 62104 2076
rect 62160 2020 62188 2076
rect 61836 1996 62188 2020
rect 61384 1964 61436 1970
rect 61384 1906 61436 1912
rect 61836 1940 61864 1996
rect 61920 1940 61944 1996
rect 62000 1940 62024 1996
rect 62080 1940 62104 1996
rect 62160 1940 62188 1996
rect 61108 1896 61160 1902
rect 61108 1838 61160 1844
rect 61016 1556 61068 1562
rect 61016 1498 61068 1504
rect 61120 800 61148 1838
rect 61836 1658 62188 1940
rect 61836 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 62188 1658
rect 61836 1040 62188 1606
rect 62316 1306 62344 2382
rect 62948 2304 63000 2310
rect 62948 2246 63000 2252
rect 62960 1970 62988 2246
rect 62948 1964 63000 1970
rect 62948 1906 63000 1912
rect 62396 1760 62448 1766
rect 62396 1702 62448 1708
rect 62408 1358 62436 1702
rect 62764 1420 62816 1426
rect 62764 1362 62816 1368
rect 62224 1278 62344 1306
rect 62396 1352 62448 1358
rect 62396 1294 62448 1300
rect 62224 800 62252 1278
rect 62776 800 62804 1362
rect 63052 1358 63080 2790
rect 63592 2372 63644 2378
rect 63592 2314 63644 2320
rect 63604 2106 63632 2314
rect 63696 2310 63724 6394
rect 63788 6186 63816 11834
rect 63880 6254 63908 12022
rect 63972 6322 64000 45698
rect 64188 44588 64540 54292
rect 64188 44532 64216 44588
rect 64272 44532 64296 44588
rect 64352 44532 64376 44588
rect 64432 44532 64456 44588
rect 64512 44532 64540 44588
rect 64188 44508 64540 44532
rect 64188 44452 64216 44508
rect 64272 44452 64296 44508
rect 64352 44452 64376 44508
rect 64432 44452 64456 44508
rect 64512 44452 64540 44508
rect 64188 44428 64540 44452
rect 64188 44372 64216 44428
rect 64272 44372 64296 44428
rect 64352 44372 64376 44428
rect 64432 44372 64456 44428
rect 64512 44372 64540 44428
rect 64188 44348 64540 44372
rect 64188 44292 64216 44348
rect 64272 44292 64296 44348
rect 64352 44292 64376 44348
rect 64432 44292 64456 44348
rect 64512 44292 64540 44348
rect 64052 43852 64104 43858
rect 64052 43794 64104 43800
rect 64064 11257 64092 43794
rect 64188 34588 64540 44292
rect 64188 34532 64216 34588
rect 64272 34532 64296 34588
rect 64352 34532 64376 34588
rect 64432 34532 64456 34588
rect 64512 34532 64540 34588
rect 64188 34508 64540 34532
rect 64188 34452 64216 34508
rect 64272 34452 64296 34508
rect 64352 34452 64376 34508
rect 64432 34452 64456 34508
rect 64512 34452 64540 34508
rect 64188 34428 64540 34452
rect 64188 34372 64216 34428
rect 64272 34372 64296 34428
rect 64352 34372 64376 34428
rect 64432 34372 64456 34428
rect 64512 34372 64540 34428
rect 64188 34348 64540 34372
rect 64188 34292 64216 34348
rect 64272 34292 64296 34348
rect 64352 34292 64376 34348
rect 64432 34292 64456 34348
rect 64512 34292 64540 34348
rect 64188 24588 64540 34292
rect 64188 24532 64216 24588
rect 64272 24532 64296 24588
rect 64352 24532 64376 24588
rect 64432 24532 64456 24588
rect 64512 24532 64540 24588
rect 64188 24508 64540 24532
rect 64188 24452 64216 24508
rect 64272 24452 64296 24508
rect 64352 24452 64376 24508
rect 64432 24452 64456 24508
rect 64512 24452 64540 24508
rect 64188 24428 64540 24452
rect 64188 24372 64216 24428
rect 64272 24372 64296 24428
rect 64352 24372 64376 24428
rect 64432 24372 64456 24428
rect 64512 24372 64540 24428
rect 64188 24348 64540 24372
rect 64188 24292 64216 24348
rect 64272 24292 64296 24348
rect 64352 24292 64376 24348
rect 64432 24292 64456 24348
rect 64512 24292 64540 24348
rect 64188 14588 64540 24292
rect 64188 14532 64216 14588
rect 64272 14532 64296 14588
rect 64352 14532 64376 14588
rect 64432 14532 64456 14588
rect 64512 14532 64540 14588
rect 64188 14508 64540 14532
rect 64188 14452 64216 14508
rect 64272 14452 64296 14508
rect 64352 14452 64376 14508
rect 64432 14452 64456 14508
rect 64512 14452 64540 14508
rect 64188 14428 64540 14452
rect 64188 14372 64216 14428
rect 64272 14372 64296 14428
rect 64352 14372 64376 14428
rect 64432 14372 64456 14428
rect 64512 14372 64540 14428
rect 64188 14348 64540 14372
rect 64188 14292 64216 14348
rect 64272 14292 64296 14348
rect 64352 14292 64376 14348
rect 64432 14292 64456 14348
rect 64512 14292 64540 14348
rect 64050 11248 64106 11257
rect 64050 11183 64106 11192
rect 64052 11076 64104 11082
rect 64052 11018 64104 11024
rect 64064 7993 64092 11018
rect 64050 7984 64106 7993
rect 64050 7919 64106 7928
rect 63960 6316 64012 6322
rect 63960 6258 64012 6264
rect 63868 6248 63920 6254
rect 63868 6190 63920 6196
rect 63776 6180 63828 6186
rect 63776 6122 63828 6128
rect 63776 5908 63828 5914
rect 63776 5850 63828 5856
rect 63788 5098 63816 5850
rect 64188 5466 64540 14292
rect 64616 7818 64644 67594
rect 64880 66496 64932 66502
rect 64880 66438 64932 66444
rect 64892 64326 64920 66438
rect 65432 65680 65484 65686
rect 65432 65622 65484 65628
rect 64880 64320 64932 64326
rect 64880 64262 64932 64268
rect 64892 62150 64920 64262
rect 65340 63572 65392 63578
rect 65340 63514 65392 63520
rect 64880 62144 64932 62150
rect 64880 62086 64932 62092
rect 64892 60246 64920 62086
rect 65248 61328 65300 61334
rect 65248 61270 65300 61276
rect 64880 60240 64932 60246
rect 64880 60182 64932 60188
rect 64892 58070 64920 60182
rect 65156 59152 65208 59158
rect 65156 59094 65208 59100
rect 64880 58064 64932 58070
rect 64880 58006 64932 58012
rect 64892 55622 64920 58006
rect 64880 55616 64932 55622
rect 64880 55558 64932 55564
rect 64892 53582 64920 55558
rect 64880 53576 64932 53582
rect 64880 53518 64932 53524
rect 64892 51542 64920 53518
rect 64880 51536 64932 51542
rect 64880 51478 64932 51484
rect 64788 47048 64840 47054
rect 64788 46990 64840 46996
rect 64696 33992 64748 33998
rect 64696 33934 64748 33940
rect 64604 7812 64656 7818
rect 64604 7754 64656 7760
rect 64604 7132 64656 7138
rect 64604 7074 64656 7080
rect 64616 6186 64644 7074
rect 64708 6526 64736 33934
rect 64696 6520 64748 6526
rect 64696 6462 64748 6468
rect 64696 6248 64748 6254
rect 64696 6190 64748 6196
rect 64604 6180 64656 6186
rect 64604 6122 64656 6128
rect 64188 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64540 5466
rect 63776 5092 63828 5098
rect 63776 5034 63828 5040
rect 64188 4588 64540 5414
rect 64188 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64540 4588
rect 64188 4508 64540 4532
rect 64188 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64540 4508
rect 64188 4428 64540 4452
rect 64188 4378 64216 4428
rect 64272 4378 64296 4428
rect 64352 4378 64376 4428
rect 64432 4378 64456 4428
rect 64512 4378 64540 4428
rect 64188 4326 64210 4378
rect 64272 4372 64274 4378
rect 64454 4372 64456 4378
rect 64262 4348 64274 4372
rect 64326 4348 64338 4372
rect 64390 4348 64402 4372
rect 64454 4348 64466 4372
rect 64272 4326 64274 4348
rect 64454 4326 64456 4348
rect 64518 4326 64540 4378
rect 64188 4292 64216 4326
rect 64272 4292 64296 4326
rect 64352 4292 64376 4326
rect 64432 4292 64456 4326
rect 64512 4292 64540 4326
rect 64188 3290 64540 4292
rect 64188 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64540 3290
rect 63684 2304 63736 2310
rect 63684 2246 63736 2252
rect 64188 2202 64540 3238
rect 64708 3126 64736 6190
rect 64800 5953 64828 46990
rect 64880 44872 64932 44878
rect 64880 44814 64932 44820
rect 64892 35894 64920 44814
rect 65064 41744 65116 41750
rect 65064 41686 65116 41692
rect 64972 40996 65024 41002
rect 64972 40938 65024 40944
rect 64984 40905 65012 40938
rect 64970 40896 65026 40905
rect 64970 40831 65026 40840
rect 65076 39846 65104 41686
rect 65064 39840 65116 39846
rect 65064 39782 65116 39788
rect 64972 38888 65024 38894
rect 64970 38856 64972 38865
rect 65024 38856 65026 38865
rect 64970 38791 65026 38800
rect 65076 37398 65104 39782
rect 65064 37392 65116 37398
rect 65064 37334 65116 37340
rect 64892 35866 65012 35894
rect 64880 35216 64932 35222
rect 64880 35158 64932 35164
rect 64892 33318 64920 35158
rect 64880 33312 64932 33318
rect 64880 33254 64932 33260
rect 64892 31142 64920 33254
rect 64880 31136 64932 31142
rect 64880 31078 64932 31084
rect 64892 28694 64920 31078
rect 64880 28688 64932 28694
rect 64880 28630 64932 28636
rect 64892 27130 64920 28630
rect 64880 27124 64932 27130
rect 64880 27066 64932 27072
rect 64984 23866 65012 35866
rect 65076 35222 65104 37334
rect 65064 35216 65116 35222
rect 65064 35158 65116 35164
rect 65168 30938 65196 59094
rect 65260 32450 65288 61270
rect 65352 33114 65380 63514
rect 65444 33658 65472 65622
rect 65536 36378 65564 69974
rect 65892 67856 65944 67862
rect 65892 67798 65944 67804
rect 65708 65408 65760 65414
rect 65708 65350 65760 65356
rect 65616 52488 65668 52494
rect 65616 52430 65668 52436
rect 65628 52154 65656 52430
rect 65616 52148 65668 52154
rect 65616 52090 65668 52096
rect 65524 36372 65576 36378
rect 65524 36314 65576 36320
rect 65522 34776 65578 34785
rect 65522 34711 65578 34720
rect 65536 34610 65564 34711
rect 65524 34604 65576 34610
rect 65524 34546 65576 34552
rect 65616 33924 65668 33930
rect 65616 33866 65668 33872
rect 65432 33652 65484 33658
rect 65432 33594 65484 33600
rect 65628 33289 65656 33866
rect 65614 33280 65670 33289
rect 65614 33215 65670 33224
rect 65340 33108 65392 33114
rect 65340 33050 65392 33056
rect 65260 32422 65380 32450
rect 65248 32224 65300 32230
rect 65248 32166 65300 32172
rect 65156 30932 65208 30938
rect 65156 30874 65208 30880
rect 65156 24336 65208 24342
rect 65156 24278 65208 24284
rect 64972 23860 65024 23866
rect 64972 23802 65024 23808
rect 65168 22166 65196 24278
rect 65156 22160 65208 22166
rect 65156 22102 65208 22108
rect 65168 20262 65196 22102
rect 65156 20256 65208 20262
rect 65156 20198 65208 20204
rect 65064 19168 65116 19174
rect 65064 19110 65116 19116
rect 64972 14816 65024 14822
rect 64972 14758 65024 14764
rect 64880 12776 64932 12782
rect 64878 12744 64880 12753
rect 64932 12744 64934 12753
rect 64878 12679 64934 12688
rect 64878 12608 64934 12617
rect 64878 12543 64934 12552
rect 64892 11801 64920 12543
rect 64878 11792 64934 11801
rect 64878 11727 64934 11736
rect 64880 10464 64932 10470
rect 64880 10406 64932 10412
rect 64892 6866 64920 10406
rect 64984 7750 65012 14758
rect 64972 7744 65024 7750
rect 64972 7686 65024 7692
rect 65076 7614 65104 19110
rect 65168 18018 65196 20198
rect 65156 18012 65208 18018
rect 65156 17954 65208 17960
rect 65168 15638 65196 17954
rect 65156 15632 65208 15638
rect 65156 15574 65208 15580
rect 65168 13734 65196 15574
rect 65156 13728 65208 13734
rect 65156 13670 65208 13676
rect 65168 11286 65196 13670
rect 65156 11280 65208 11286
rect 65156 11222 65208 11228
rect 65168 9382 65196 11222
rect 65156 9376 65208 9382
rect 65156 9318 65208 9324
rect 65064 7608 65116 7614
rect 65064 7550 65116 7556
rect 65064 7064 65116 7070
rect 65064 7006 65116 7012
rect 64880 6860 64932 6866
rect 64880 6802 64932 6808
rect 64972 6792 65024 6798
rect 64972 6734 65024 6740
rect 64984 6594 65012 6734
rect 65076 6662 65104 7006
rect 65064 6656 65116 6662
rect 65064 6598 65116 6604
rect 64972 6588 65024 6594
rect 64972 6530 65024 6536
rect 64878 6352 64934 6361
rect 64878 6287 64934 6296
rect 64972 6316 65024 6322
rect 64786 5944 64842 5953
rect 64786 5879 64842 5888
rect 64788 5568 64840 5574
rect 64788 5510 64840 5516
rect 64696 3120 64748 3126
rect 64696 3062 64748 3068
rect 64800 3058 64828 5510
rect 64892 3097 64920 6287
rect 64972 6258 65024 6264
rect 64984 5545 65012 6258
rect 64970 5536 65026 5545
rect 64970 5471 65026 5480
rect 65168 4758 65196 9318
rect 65260 5914 65288 32166
rect 65352 32026 65380 32422
rect 65340 32020 65392 32026
rect 65340 31962 65392 31968
rect 65340 30048 65392 30054
rect 65340 29990 65392 29996
rect 65248 5908 65300 5914
rect 65248 5850 65300 5856
rect 65352 5642 65380 29990
rect 65432 25696 65484 25702
rect 65432 25638 65484 25644
rect 65340 5636 65392 5642
rect 65340 5578 65392 5584
rect 65444 5166 65472 25638
rect 65524 23520 65576 23526
rect 65524 23462 65576 23468
rect 65432 5160 65484 5166
rect 65432 5102 65484 5108
rect 65156 4752 65208 4758
rect 65156 4694 65208 4700
rect 65536 4214 65564 23462
rect 65616 16992 65668 16998
rect 65616 16934 65668 16940
rect 65628 7886 65656 16934
rect 65616 7880 65668 7886
rect 65616 7822 65668 7828
rect 65720 7342 65748 65350
rect 65800 56704 65852 56710
rect 65800 56646 65852 56652
rect 65708 7336 65760 7342
rect 65708 7278 65760 7284
rect 65812 7274 65840 56646
rect 65904 35290 65932 67798
rect 65892 35284 65944 35290
rect 65892 35226 65944 35232
rect 65892 27872 65944 27878
rect 65892 27814 65944 27820
rect 65800 7268 65852 7274
rect 65800 7210 65852 7216
rect 65904 7206 65932 27814
rect 65892 7200 65944 7206
rect 65892 7142 65944 7148
rect 65800 6860 65852 6866
rect 65800 6802 65852 6808
rect 65708 6724 65760 6730
rect 65708 6666 65760 6672
rect 65524 4208 65576 4214
rect 65524 4150 65576 4156
rect 64878 3088 64934 3097
rect 64788 3052 64840 3058
rect 64878 3023 64934 3032
rect 64788 2994 64840 3000
rect 64604 2848 64656 2854
rect 64604 2790 64656 2796
rect 64188 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64540 2202
rect 63592 2100 63644 2106
rect 63592 2042 63644 2048
rect 63868 1896 63920 1902
rect 63868 1838 63920 1844
rect 63880 1562 63908 1838
rect 63868 1556 63920 1562
rect 63868 1498 63920 1504
rect 63040 1352 63092 1358
rect 63040 1294 63092 1300
rect 63868 1352 63920 1358
rect 63868 1294 63920 1300
rect 63880 800 63908 1294
rect 64188 1114 64540 2150
rect 64616 1970 64644 2790
rect 65720 2514 65748 6666
rect 65708 2508 65760 2514
rect 65708 2450 65760 2456
rect 65524 2440 65576 2446
rect 65524 2382 65576 2388
rect 64604 1964 64656 1970
rect 64604 1906 64656 1912
rect 64696 1896 64748 1902
rect 64696 1838 64748 1844
rect 64188 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64540 1114
rect 64188 1040 64540 1062
rect 64432 870 64552 898
rect 64432 800 64460 870
rect 44652 734 44864 762
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64524 762 64552 870
rect 64708 762 64736 1838
rect 65156 1760 65208 1766
rect 65156 1702 65208 1708
rect 65168 1358 65196 1702
rect 65156 1352 65208 1358
rect 65156 1294 65208 1300
rect 65536 800 65564 2382
rect 65812 1834 65840 6802
rect 65996 5778 66024 71878
rect 66076 36576 66128 36582
rect 66076 36518 66128 36524
rect 66088 6497 66116 36518
rect 66074 6488 66130 6497
rect 66074 6423 66130 6432
rect 66180 5778 66208 74054
rect 66272 39642 66300 76502
rect 66352 72208 66404 72214
rect 66352 72150 66404 72156
rect 66260 39636 66312 39642
rect 66260 39578 66312 39584
rect 66364 37194 66392 72150
rect 66456 40730 66484 78678
rect 66536 69012 66588 69018
rect 66536 68954 66588 68960
rect 66444 40724 66496 40730
rect 66444 40666 66496 40672
rect 66352 37188 66404 37194
rect 66352 37130 66404 37136
rect 66352 36168 66404 36174
rect 66352 36110 66404 36116
rect 66260 31816 66312 31822
rect 66260 31758 66312 31764
rect 66272 6458 66300 31758
rect 66260 6452 66312 6458
rect 66260 6394 66312 6400
rect 66364 6236 66392 36110
rect 66548 35766 66576 68954
rect 66904 53168 66956 53174
rect 66904 53110 66956 53116
rect 66628 51536 66680 51542
rect 66628 51478 66680 51484
rect 66536 35760 66588 35766
rect 66536 35702 66588 35708
rect 66444 32904 66496 32910
rect 66444 32846 66496 32852
rect 66456 26234 66484 32846
rect 66536 30728 66588 30734
rect 66536 30670 66588 30676
rect 66548 26874 66576 30670
rect 66640 27062 66668 51478
rect 66812 46980 66864 46986
rect 66812 46922 66864 46928
rect 66720 33448 66772 33454
rect 66720 33390 66772 33396
rect 66628 27056 66680 27062
rect 66628 26998 66680 27004
rect 66548 26846 66668 26874
rect 66456 26206 66576 26234
rect 66444 24200 66496 24206
rect 66444 24142 66496 24148
rect 66456 23497 66484 24142
rect 66442 23488 66498 23497
rect 66442 23423 66498 23432
rect 66444 23112 66496 23118
rect 66444 23054 66496 23060
rect 66456 22409 66484 23054
rect 66442 22400 66498 22409
rect 66442 22335 66498 22344
rect 66444 22228 66496 22234
rect 66444 22170 66496 22176
rect 66272 6208 66392 6236
rect 65984 5772 66036 5778
rect 65984 5714 66036 5720
rect 66168 5772 66220 5778
rect 66168 5714 66220 5720
rect 66272 5658 66300 6208
rect 66456 5658 66484 22170
rect 66180 5630 66300 5658
rect 66364 5630 66484 5658
rect 66180 2582 66208 5630
rect 66364 3602 66392 5630
rect 66444 5568 66496 5574
rect 66444 5510 66496 5516
rect 66352 3596 66404 3602
rect 66352 3538 66404 3544
rect 66456 3058 66484 5510
rect 66548 4078 66576 26206
rect 66640 4146 66668 26846
rect 66732 6866 66760 33390
rect 66824 11082 66852 46922
rect 66916 34202 66944 53110
rect 67008 42770 67036 83098
rect 69664 83020 69716 83026
rect 69664 82962 69716 82968
rect 67088 80980 67140 80986
rect 67088 80922 67140 80928
rect 66996 42764 67048 42770
rect 66996 42706 67048 42712
rect 67100 41818 67128 80922
rect 68468 76492 68520 76498
rect 68468 76434 68520 76440
rect 67640 74656 67692 74662
rect 67640 74598 67692 74604
rect 67548 54800 67600 54806
rect 67548 54742 67600 54748
rect 67364 50448 67416 50454
rect 67364 50390 67416 50396
rect 67180 47048 67232 47054
rect 67180 46990 67232 46996
rect 67088 41812 67140 41818
rect 67088 41754 67140 41760
rect 66996 38344 67048 38350
rect 66996 38286 67048 38292
rect 66904 34196 66956 34202
rect 66904 34138 66956 34144
rect 67008 31090 67036 38286
rect 67088 35080 67140 35086
rect 67088 35022 67140 35028
rect 66916 31062 67036 31090
rect 66812 11076 66864 11082
rect 66812 11018 66864 11024
rect 66720 6860 66772 6866
rect 66720 6802 66772 6808
rect 66628 4140 66680 4146
rect 66628 4082 66680 4088
rect 66536 4072 66588 4078
rect 66536 4014 66588 4020
rect 66444 3052 66496 3058
rect 66444 2994 66496 3000
rect 66260 2848 66312 2854
rect 66260 2790 66312 2796
rect 66168 2576 66220 2582
rect 66168 2518 66220 2524
rect 66076 2304 66128 2310
rect 66076 2246 66128 2252
rect 66088 1970 66116 2246
rect 66076 1964 66128 1970
rect 66076 1906 66128 1912
rect 65800 1828 65852 1834
rect 65800 1770 65852 1776
rect 66272 1358 66300 2790
rect 66916 2038 66944 31062
rect 66996 29640 67048 29646
rect 66996 29582 67048 29588
rect 67008 6254 67036 29582
rect 67100 6730 67128 35022
rect 67192 7449 67220 46990
rect 67272 37256 67324 37262
rect 67272 37198 67324 37204
rect 67178 7440 67234 7449
rect 67178 7375 67234 7384
rect 67088 6724 67140 6730
rect 67088 6666 67140 6672
rect 66996 6248 67048 6254
rect 66996 6190 67048 6196
rect 67284 2530 67312 37198
rect 67376 28694 67404 50390
rect 67456 39432 67508 39438
rect 67456 39374 67508 39380
rect 67364 28688 67416 28694
rect 67364 28630 67416 28636
rect 67364 28552 67416 28558
rect 67364 28494 67416 28500
rect 67376 26489 67404 28494
rect 67362 26480 67418 26489
rect 67362 26415 67418 26424
rect 67364 26376 67416 26382
rect 67364 26318 67416 26324
rect 67376 3534 67404 26318
rect 67364 3528 67416 3534
rect 67364 3470 67416 3476
rect 67284 2502 67404 2530
rect 67468 2514 67496 39374
rect 67560 28762 67588 54742
rect 67652 38554 67680 74598
rect 68100 57044 68152 57050
rect 68100 56986 68152 56992
rect 67732 44464 67784 44470
rect 67732 44406 67784 44412
rect 67640 38548 67692 38554
rect 67640 38490 67692 38496
rect 67548 28756 67600 28762
rect 67548 28698 67600 28704
rect 67548 28620 67600 28626
rect 67548 28562 67600 28568
rect 67560 27554 67588 28562
rect 67560 27526 67680 27554
rect 67548 27464 67600 27470
rect 67548 27406 67600 27412
rect 67560 26194 67588 27406
rect 67652 26586 67680 27526
rect 67640 26580 67692 26586
rect 67640 26522 67692 26528
rect 67560 26166 67680 26194
rect 67546 26072 67602 26081
rect 67546 26007 67602 26016
rect 67272 2440 67324 2446
rect 67272 2382 67324 2388
rect 67284 2106 67312 2382
rect 67272 2100 67324 2106
rect 67272 2042 67324 2048
rect 66904 2032 66956 2038
rect 66904 1974 66956 1980
rect 67180 1964 67232 1970
rect 67180 1906 67232 1912
rect 66260 1352 66312 1358
rect 66260 1294 66312 1300
rect 66076 1284 66128 1290
rect 66076 1226 66128 1232
rect 66088 800 66116 1226
rect 67192 800 67220 1906
rect 67376 1222 67404 2502
rect 67456 2508 67508 2514
rect 67456 2450 67508 2456
rect 67560 2378 67588 26007
rect 67652 23746 67680 26166
rect 67744 24410 67772 44406
rect 67916 40928 67968 40934
rect 67916 40870 67968 40876
rect 67732 24404 67784 24410
rect 67732 24346 67784 24352
rect 67652 23718 67772 23746
rect 67640 23656 67692 23662
rect 67638 23624 67640 23633
rect 67692 23624 67694 23633
rect 67638 23559 67694 23568
rect 67744 22234 67772 23718
rect 67732 22228 67784 22234
rect 67732 22170 67784 22176
rect 67824 18964 67876 18970
rect 67824 18906 67876 18912
rect 67640 14612 67692 14618
rect 67640 14554 67692 14560
rect 67652 5846 67680 14554
rect 67732 12640 67784 12646
rect 67732 12582 67784 12588
rect 67744 6390 67772 12582
rect 67836 7546 67864 18906
rect 67824 7540 67876 7546
rect 67824 7482 67876 7488
rect 67928 6798 67956 40870
rect 68008 38752 68060 38758
rect 68008 38694 68060 38700
rect 67916 6792 67968 6798
rect 67916 6734 67968 6740
rect 67732 6384 67784 6390
rect 67732 6326 67784 6332
rect 67640 5840 67692 5846
rect 67640 5782 67692 5788
rect 68020 4486 68048 38694
rect 68112 29850 68140 56986
rect 68192 52692 68244 52698
rect 68192 52634 68244 52640
rect 68100 29844 68152 29850
rect 68100 29786 68152 29792
rect 68204 27606 68232 52634
rect 68376 46028 68428 46034
rect 68376 45970 68428 45976
rect 68284 44532 68336 44538
rect 68284 44474 68336 44480
rect 68192 27600 68244 27606
rect 68192 27542 68244 27548
rect 68100 27124 68152 27130
rect 68100 27066 68152 27072
rect 68112 7478 68140 27066
rect 68296 23322 68324 44474
rect 68284 23316 68336 23322
rect 68284 23258 68336 23264
rect 68192 21140 68244 21146
rect 68192 21082 68244 21088
rect 68100 7472 68152 7478
rect 68100 7414 68152 7420
rect 68204 6118 68232 21082
rect 68388 6186 68416 45970
rect 68376 6180 68428 6186
rect 68376 6122 68428 6128
rect 68192 6112 68244 6118
rect 68192 6054 68244 6060
rect 68480 5778 68508 76434
rect 69020 63436 69072 63442
rect 69020 63378 69072 63384
rect 68560 47524 68612 47530
rect 68560 47466 68612 47472
rect 68468 5772 68520 5778
rect 68468 5714 68520 5720
rect 68100 5568 68152 5574
rect 68100 5510 68152 5516
rect 68008 4480 68060 4486
rect 68008 4422 68060 4428
rect 68112 3058 68140 5510
rect 68572 4622 68600 47466
rect 68744 43104 68796 43110
rect 68744 43046 68796 43052
rect 68652 25492 68704 25498
rect 68652 25434 68704 25440
rect 68664 6322 68692 25434
rect 68652 6316 68704 6322
rect 68652 6258 68704 6264
rect 68756 4826 68784 43046
rect 68836 23248 68888 23254
rect 68836 23190 68888 23196
rect 68848 6662 68876 23190
rect 68836 6656 68888 6662
rect 68836 6598 68888 6604
rect 69032 5817 69060 63378
rect 69112 54664 69164 54670
rect 69112 54606 69164 54612
rect 69018 5808 69074 5817
rect 69018 5743 69074 5752
rect 69124 5409 69152 54606
rect 69204 40520 69256 40526
rect 69204 40462 69256 40468
rect 69110 5400 69166 5409
rect 69110 5335 69166 5344
rect 68744 4820 68796 4826
rect 68744 4762 68796 4768
rect 68560 4616 68612 4622
rect 68560 4558 68612 4564
rect 68100 3052 68152 3058
rect 68100 2994 68152 3000
rect 68284 2848 68336 2854
rect 68284 2790 68336 2796
rect 67548 2372 67600 2378
rect 67548 2314 67600 2320
rect 67732 1420 67784 1426
rect 67732 1362 67784 1368
rect 67364 1216 67416 1222
rect 67364 1158 67416 1164
rect 67744 800 67772 1362
rect 68296 1358 68324 2790
rect 69216 2038 69244 40462
rect 69296 36304 69348 36310
rect 69296 36246 69348 36252
rect 69308 4554 69336 36246
rect 69388 21548 69440 21554
rect 69388 21490 69440 21496
rect 69400 6866 69428 21490
rect 69388 6860 69440 6866
rect 69388 6802 69440 6808
rect 69676 5302 69704 82962
rect 71836 82236 72188 83206
rect 71836 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 72188 82236
rect 71836 82170 72188 82180
rect 71836 82118 71858 82170
rect 71910 82156 71922 82170
rect 71974 82156 71986 82170
rect 72038 82156 72050 82170
rect 72102 82156 72114 82170
rect 71920 82118 71922 82156
rect 72102 82118 72104 82156
rect 72166 82118 72188 82170
rect 71836 82100 71864 82118
rect 71920 82100 71944 82118
rect 72000 82100 72024 82118
rect 72080 82100 72104 82118
rect 72160 82100 72188 82118
rect 71836 82076 72188 82100
rect 71836 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 72188 82076
rect 71836 81996 72188 82020
rect 71836 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 72188 81996
rect 71836 81082 72188 81940
rect 71836 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 72188 81082
rect 69756 80844 69808 80850
rect 69756 80786 69808 80792
rect 69664 5296 69716 5302
rect 69664 5238 69716 5244
rect 69768 5098 69796 80786
rect 71836 79994 72188 81030
rect 71836 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 72188 79994
rect 71836 78906 72188 79942
rect 71836 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 72188 78906
rect 69940 78668 69992 78674
rect 69940 78610 69992 78616
rect 69952 5166 69980 78610
rect 71836 77818 72188 78854
rect 71836 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 72188 77818
rect 71836 76730 72188 77766
rect 71836 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 72188 76730
rect 71836 75642 72188 76678
rect 71836 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 72188 75642
rect 71836 74554 72188 75590
rect 71836 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 72188 74554
rect 71836 73466 72188 74502
rect 71836 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 72188 73466
rect 71836 72378 72188 73414
rect 71836 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 72188 72378
rect 71836 72236 72188 72326
rect 71836 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 72188 72236
rect 71836 72156 72188 72180
rect 71836 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 72188 72156
rect 71836 72076 72188 72100
rect 71836 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 72188 72076
rect 71836 71996 72188 72020
rect 71836 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 72188 71996
rect 71836 71290 72188 71940
rect 71836 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 72188 71290
rect 71836 70202 72188 71238
rect 71836 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 72188 70202
rect 71836 69114 72188 70150
rect 71836 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 72188 69114
rect 71836 68026 72188 69062
rect 71836 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 72188 68026
rect 71836 66938 72188 67974
rect 71836 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 72188 66938
rect 71836 65850 72188 66886
rect 71836 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 72188 65850
rect 71836 64762 72188 65798
rect 71836 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 72188 64762
rect 71836 63674 72188 64710
rect 71836 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 72188 63674
rect 71836 62586 72188 63622
rect 71836 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 72188 62586
rect 71836 62236 72188 62534
rect 71836 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 72188 62236
rect 71836 62156 72188 62180
rect 71836 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 72188 62156
rect 71836 62076 72188 62100
rect 71836 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 72188 62076
rect 71836 61996 72188 62020
rect 71836 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 72188 61996
rect 71836 61498 72188 61940
rect 71836 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 72188 61498
rect 71836 60410 72188 61446
rect 71836 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 72188 60410
rect 71836 59322 72188 60358
rect 71836 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 72188 59322
rect 70768 59084 70820 59090
rect 70768 59026 70820 59032
rect 70492 43308 70544 43314
rect 70492 43250 70544 43256
rect 70032 42696 70084 42702
rect 70032 42638 70084 42644
rect 69940 5160 69992 5166
rect 69940 5102 69992 5108
rect 69756 5092 69808 5098
rect 69756 5034 69808 5040
rect 69848 5024 69900 5030
rect 69848 4966 69900 4972
rect 69296 4548 69348 4554
rect 69296 4490 69348 4496
rect 69860 3058 69888 4966
rect 69848 3052 69900 3058
rect 69848 2994 69900 3000
rect 69664 2848 69716 2854
rect 69664 2790 69716 2796
rect 69388 2304 69440 2310
rect 69388 2246 69440 2252
rect 69204 2032 69256 2038
rect 69204 1974 69256 1980
rect 69400 1970 69428 2246
rect 69676 1970 69704 2790
rect 69940 2440 69992 2446
rect 69940 2382 69992 2388
rect 69388 1964 69440 1970
rect 69388 1906 69440 1912
rect 69664 1964 69716 1970
rect 69664 1906 69716 1912
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 68284 1352 68336 1358
rect 68284 1294 68336 1300
rect 68836 1352 68888 1358
rect 68836 1294 68888 1300
rect 68848 800 68876 1294
rect 69400 800 69428 1770
rect 69952 1562 69980 2382
rect 69940 1556 69992 1562
rect 69940 1498 69992 1504
rect 70044 1290 70072 42638
rect 70124 41608 70176 41614
rect 70124 41550 70176 41556
rect 70136 2038 70164 41550
rect 70504 5273 70532 43250
rect 70584 35692 70636 35698
rect 70584 35634 70636 35640
rect 70490 5264 70546 5273
rect 70490 5199 70546 5208
rect 70492 2440 70544 2446
rect 70492 2382 70544 2388
rect 70124 2032 70176 2038
rect 70124 1974 70176 1980
rect 70032 1284 70084 1290
rect 70032 1226 70084 1232
rect 70504 800 70532 2382
rect 70596 2106 70624 35634
rect 70676 26988 70728 26994
rect 70676 26930 70728 26936
rect 70688 2650 70716 26930
rect 70780 4690 70808 59026
rect 71836 58234 72188 59270
rect 71836 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 72188 58234
rect 71836 57146 72188 58182
rect 71836 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 72188 57146
rect 71836 56058 72188 57094
rect 71836 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 72188 56058
rect 71836 54970 72188 56006
rect 71836 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 72188 54970
rect 71836 53882 72188 54918
rect 71836 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 72188 53882
rect 71836 52794 72188 53830
rect 71836 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 72188 52794
rect 71836 52236 72188 52742
rect 71836 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 72188 52236
rect 71836 52156 72188 52180
rect 71836 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 72188 52156
rect 71836 52076 72188 52100
rect 71836 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 72188 52076
rect 71836 51996 72188 52020
rect 71836 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 72188 51996
rect 71836 51706 72188 51940
rect 71836 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 72188 51706
rect 71836 50618 72188 51654
rect 71836 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 72188 50618
rect 71836 49530 72188 50566
rect 71836 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 72188 49530
rect 71836 48442 72188 49478
rect 71836 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 72188 48442
rect 71836 47354 72188 48390
rect 71836 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 72188 47354
rect 71836 46266 72188 47302
rect 71836 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 72188 46266
rect 71836 45178 72188 46214
rect 71836 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 72188 45178
rect 71836 44090 72188 45126
rect 71836 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 72188 44090
rect 71836 43002 72188 44038
rect 71836 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 72188 43002
rect 71836 42236 72188 42950
rect 71836 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 72188 42236
rect 71836 42156 72188 42180
rect 71836 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 72188 42156
rect 71836 42076 72188 42100
rect 71836 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 72188 42076
rect 71836 41996 72188 42020
rect 71836 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 72188 41996
rect 71836 41914 72188 41940
rect 71836 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 72188 41914
rect 71836 40826 72188 41862
rect 71836 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 72188 40826
rect 71836 39738 72188 40774
rect 71836 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 72188 39738
rect 71836 38650 72188 39686
rect 71836 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 72188 38650
rect 71836 37562 72188 38598
rect 71836 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 72188 37562
rect 71836 36474 72188 37510
rect 71836 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 72188 36474
rect 71836 35386 72188 36422
rect 71836 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 72188 35386
rect 71836 34298 72188 35334
rect 71836 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 72188 34298
rect 71836 33210 72188 34246
rect 71836 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 72188 33210
rect 71836 32236 72188 33158
rect 71836 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 72188 32236
rect 71836 32156 72188 32180
rect 71836 32122 71864 32156
rect 71920 32122 71944 32156
rect 72000 32122 72024 32156
rect 72080 32122 72104 32156
rect 72160 32122 72188 32156
rect 71836 32070 71858 32122
rect 71920 32100 71922 32122
rect 72102 32100 72104 32122
rect 71910 32076 71922 32100
rect 71974 32076 71986 32100
rect 72038 32076 72050 32100
rect 72102 32076 72114 32100
rect 71920 32070 71922 32076
rect 72102 32070 72104 32076
rect 72166 32070 72188 32122
rect 71836 32020 71864 32070
rect 71920 32020 71944 32070
rect 72000 32020 72024 32070
rect 72080 32020 72104 32070
rect 72160 32020 72188 32070
rect 71836 31996 72188 32020
rect 71836 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 72188 31996
rect 71836 31034 72188 31940
rect 71836 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 72188 31034
rect 71836 29946 72188 30982
rect 71836 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 72188 29946
rect 71836 28858 72188 29894
rect 71836 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 72188 28858
rect 71836 27770 72188 28806
rect 71836 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 72188 27770
rect 71836 26682 72188 27718
rect 71836 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 72188 26682
rect 71836 25594 72188 26630
rect 71836 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 72188 25594
rect 71836 24506 72188 25542
rect 71836 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 72188 24506
rect 71836 23418 72188 24454
rect 71836 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 72188 23418
rect 71836 22330 72188 23366
rect 71836 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 72188 22330
rect 71836 22236 72188 22278
rect 71836 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 72188 22236
rect 71836 22156 72188 22180
rect 71836 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 72188 22156
rect 71836 22076 72188 22100
rect 71836 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 72188 22076
rect 71836 21996 72188 22020
rect 71836 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 72188 21996
rect 71836 21242 72188 21940
rect 71836 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 72188 21242
rect 71836 20154 72188 21190
rect 71836 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 72188 20154
rect 71836 19066 72188 20102
rect 71836 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 72188 19066
rect 71836 17978 72188 19014
rect 71836 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 72188 17978
rect 71836 16890 72188 17926
rect 71836 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 72188 16890
rect 71836 15802 72188 16838
rect 71836 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 72188 15802
rect 71836 14714 72188 15750
rect 71836 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 72188 14714
rect 71836 13626 72188 14662
rect 71836 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 72188 13626
rect 71836 12538 72188 13574
rect 71836 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 72188 12538
rect 71836 12236 72188 12486
rect 71836 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 72188 12236
rect 71836 12156 72188 12180
rect 71836 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 72188 12156
rect 71836 12076 72188 12100
rect 71836 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 72188 12076
rect 71836 11996 72188 12020
rect 71836 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 72188 11996
rect 71836 11450 72188 11940
rect 71836 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 72188 11450
rect 71836 10362 72188 11398
rect 71836 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 72188 10362
rect 71836 9274 72188 10310
rect 71836 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 72188 9274
rect 71836 8186 72188 9222
rect 71836 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 72188 8186
rect 71836 7098 72188 8134
rect 71836 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 72188 7098
rect 71836 6010 72188 7046
rect 71836 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 72188 6010
rect 71412 5024 71464 5030
rect 71412 4966 71464 4972
rect 70768 4684 70820 4690
rect 70768 4626 70820 4632
rect 71424 3058 71452 4966
rect 71836 4922 72188 5958
rect 74188 85978 74540 86000
rect 74188 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74540 85978
rect 74188 84890 74540 85926
rect 74188 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74540 84890
rect 74188 84588 74540 84838
rect 74188 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 74540 84588
rect 74188 84508 74540 84532
rect 74188 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 74540 84508
rect 74188 84428 74540 84452
rect 74188 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 74540 84428
rect 74188 84348 74540 84372
rect 74188 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 74540 84348
rect 74188 83802 74540 84292
rect 74188 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74540 83802
rect 74188 82714 74540 83750
rect 74188 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74540 82714
rect 74188 81626 74540 82662
rect 74188 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74540 81626
rect 74188 80538 74540 81574
rect 74188 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74540 80538
rect 74188 79450 74540 80486
rect 74188 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74540 79450
rect 74188 78362 74540 79398
rect 74188 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74540 78362
rect 74188 77274 74540 78310
rect 74188 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74540 77274
rect 74188 76186 74540 77222
rect 74188 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74540 76186
rect 74188 75098 74540 76134
rect 74188 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74540 75098
rect 74188 74588 74540 75046
rect 74188 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 74540 74588
rect 74188 74508 74540 74532
rect 74188 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 74540 74508
rect 74188 74428 74540 74452
rect 74188 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 74540 74428
rect 74188 74348 74540 74372
rect 74188 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 74540 74348
rect 74188 74010 74540 74292
rect 74188 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74540 74010
rect 74188 72922 74540 73958
rect 74188 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74540 72922
rect 74188 71834 74540 72870
rect 74188 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74540 71834
rect 74188 70746 74540 71782
rect 74188 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74540 70746
rect 74188 69658 74540 70694
rect 74188 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74540 69658
rect 74188 68570 74540 69606
rect 74188 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74540 68570
rect 74188 67482 74540 68518
rect 74188 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74540 67482
rect 74188 66394 74540 67430
rect 74188 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74540 66394
rect 74188 65306 74540 66342
rect 74188 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74540 65306
rect 74188 64588 74540 65254
rect 74188 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 74540 64588
rect 74188 64508 74540 64532
rect 74188 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 74540 64508
rect 74188 64428 74540 64452
rect 74188 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 74540 64428
rect 74188 64348 74540 64372
rect 74188 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 74540 64348
rect 74188 64218 74540 64292
rect 74188 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74540 64218
rect 74188 63130 74540 64166
rect 74188 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74540 63130
rect 74188 62042 74540 63078
rect 74188 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74540 62042
rect 74188 60954 74540 61990
rect 74188 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74540 60954
rect 74188 59866 74540 60902
rect 74188 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74540 59866
rect 74188 58778 74540 59814
rect 74188 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74540 58778
rect 74188 57690 74540 58726
rect 74188 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74540 57690
rect 74188 56602 74540 57638
rect 74188 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74540 56602
rect 74188 55514 74540 56550
rect 74188 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74540 55514
rect 74188 54588 74540 55462
rect 74188 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 74540 54588
rect 74188 54508 74540 54532
rect 74188 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 74540 54508
rect 74188 54428 74540 54452
rect 74188 54426 74216 54428
rect 74272 54426 74296 54428
rect 74352 54426 74376 54428
rect 74432 54426 74456 54428
rect 74512 54426 74540 54428
rect 74188 54374 74210 54426
rect 74272 54374 74274 54426
rect 74454 54374 74456 54426
rect 74518 54374 74540 54426
rect 74188 54372 74216 54374
rect 74272 54372 74296 54374
rect 74352 54372 74376 54374
rect 74432 54372 74456 54374
rect 74512 54372 74540 54374
rect 74188 54348 74540 54372
rect 74188 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 74540 54348
rect 74188 53338 74540 54292
rect 74188 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74540 53338
rect 74188 52250 74540 53286
rect 74188 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74540 52250
rect 74188 51162 74540 52198
rect 74188 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74540 51162
rect 74188 50074 74540 51110
rect 74188 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74540 50074
rect 74188 48986 74540 50022
rect 74188 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74540 48986
rect 74188 47898 74540 48934
rect 74188 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74540 47898
rect 74188 46810 74540 47846
rect 74188 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74540 46810
rect 74188 45722 74540 46758
rect 74188 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74540 45722
rect 74188 44634 74540 45670
rect 74188 44582 74210 44634
rect 74262 44588 74274 44634
rect 74326 44588 74338 44634
rect 74390 44588 74402 44634
rect 74454 44588 74466 44634
rect 74272 44582 74274 44588
rect 74454 44582 74456 44588
rect 74518 44582 74540 44634
rect 74188 44532 74216 44582
rect 74272 44532 74296 44582
rect 74352 44532 74376 44582
rect 74432 44532 74456 44582
rect 74512 44532 74540 44582
rect 74188 44508 74540 44532
rect 74188 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 74540 44508
rect 74188 44428 74540 44452
rect 74188 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 74540 44428
rect 74188 44348 74540 44372
rect 74188 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 74540 44348
rect 74188 43546 74540 44292
rect 74188 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74540 43546
rect 74188 42458 74540 43494
rect 74188 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74540 42458
rect 74188 41370 74540 42406
rect 74188 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74540 41370
rect 74188 40282 74540 41318
rect 74188 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74540 40282
rect 74188 39194 74540 40230
rect 74188 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74540 39194
rect 74188 38106 74540 39142
rect 74188 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74540 38106
rect 74188 37018 74540 38054
rect 74188 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74540 37018
rect 74188 35930 74540 36966
rect 74188 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74540 35930
rect 74188 34842 74540 35878
rect 74188 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74540 34842
rect 74188 34588 74540 34790
rect 74188 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 74540 34588
rect 74188 34508 74540 34532
rect 74188 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 74540 34508
rect 74188 34428 74540 34452
rect 74188 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 74540 34428
rect 74188 34348 74540 34372
rect 74188 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 74540 34348
rect 74188 33754 74540 34292
rect 74188 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74540 33754
rect 74188 32666 74540 33702
rect 74188 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74540 32666
rect 74188 31578 74540 32614
rect 74188 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74540 31578
rect 74188 30490 74540 31526
rect 74188 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74540 30490
rect 74188 29402 74540 30438
rect 74188 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74540 29402
rect 74188 28314 74540 29350
rect 74188 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74540 28314
rect 74188 27226 74540 28262
rect 74188 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74540 27226
rect 74188 26138 74540 27174
rect 74188 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74540 26138
rect 74188 25050 74540 26086
rect 74188 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74540 25050
rect 74188 24588 74540 24998
rect 74188 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 74540 24588
rect 74188 24508 74540 24532
rect 74188 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 74540 24508
rect 74188 24428 74540 24452
rect 74188 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 74540 24428
rect 74188 24348 74540 24372
rect 74188 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 74540 24348
rect 74188 23962 74540 24292
rect 74188 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74540 23962
rect 74188 22874 74540 23910
rect 74188 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74540 22874
rect 74188 21786 74540 22822
rect 74188 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74540 21786
rect 74188 20698 74540 21734
rect 74188 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74540 20698
rect 74188 19610 74540 20646
rect 74188 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74540 19610
rect 74188 18522 74540 19558
rect 74188 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74540 18522
rect 74188 17434 74540 18470
rect 74188 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74540 17434
rect 74188 16346 74540 17382
rect 74188 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74540 16346
rect 74188 15258 74540 16294
rect 74188 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74540 15258
rect 74188 14588 74540 15206
rect 74188 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 74540 14588
rect 74188 14508 74540 14532
rect 74188 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 74540 14508
rect 74188 14428 74540 14452
rect 74188 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 74540 14428
rect 74188 14348 74540 14372
rect 74188 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 74540 14348
rect 74188 14170 74540 14292
rect 74188 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74540 14170
rect 74188 13082 74540 14118
rect 74188 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74540 13082
rect 74188 11994 74540 13030
rect 74188 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74540 11994
rect 74188 10906 74540 11942
rect 74188 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74540 10906
rect 74188 9818 74540 10854
rect 74188 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74540 9818
rect 74188 8730 74540 9766
rect 74188 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74540 8730
rect 74188 7642 74540 8678
rect 74188 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74540 7642
rect 74188 6554 74540 7590
rect 74188 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74540 6554
rect 74188 5466 74540 6502
rect 74188 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74540 5466
rect 73252 5024 73304 5030
rect 73252 4966 73304 4972
rect 71836 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 72188 4922
rect 71836 3834 72188 4870
rect 71836 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 72188 3834
rect 71412 3052 71464 3058
rect 71412 2994 71464 3000
rect 71228 2848 71280 2854
rect 71228 2790 71280 2796
rect 70676 2644 70728 2650
rect 70676 2586 70728 2592
rect 71044 2304 71096 2310
rect 71044 2246 71096 2252
rect 70584 2100 70636 2106
rect 70584 2042 70636 2048
rect 71056 1970 71084 2246
rect 71044 1964 71096 1970
rect 71044 1906 71096 1912
rect 71044 1420 71096 1426
rect 71044 1362 71096 1368
rect 71056 800 71084 1362
rect 71240 1358 71268 2790
rect 71836 2746 72188 3782
rect 73264 3058 73292 4966
rect 74188 4588 74540 5414
rect 74188 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 74540 4588
rect 74188 4508 74540 4532
rect 74188 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 74540 4508
rect 74188 4428 74540 4452
rect 74188 4378 74216 4428
rect 74272 4378 74296 4428
rect 74352 4378 74376 4428
rect 74432 4378 74456 4428
rect 74512 4378 74540 4428
rect 74188 4326 74210 4378
rect 74272 4372 74274 4378
rect 74454 4372 74456 4378
rect 74262 4348 74274 4372
rect 74326 4348 74338 4372
rect 74390 4348 74402 4372
rect 74454 4348 74466 4372
rect 74272 4326 74274 4348
rect 74454 4326 74456 4348
rect 74518 4326 74540 4378
rect 74188 4292 74216 4326
rect 74272 4292 74296 4326
rect 74352 4292 74376 4326
rect 74432 4292 74456 4326
rect 74512 4292 74540 4326
rect 74188 3290 74540 4292
rect 74188 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74540 3290
rect 73252 3052 73304 3058
rect 73252 2994 73304 3000
rect 73252 2848 73304 2854
rect 73252 2790 73304 2796
rect 71836 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 72188 2746
rect 71836 2236 72188 2694
rect 71836 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 72188 2236
rect 71836 2156 72188 2180
rect 71836 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 72188 2156
rect 71836 2076 72188 2100
rect 71836 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 72188 2076
rect 71836 1996 72188 2020
rect 71836 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 72188 1996
rect 71836 1658 72188 1940
rect 72240 1896 72292 1902
rect 72240 1838 72292 1844
rect 71836 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 72188 1658
rect 71228 1352 71280 1358
rect 71228 1294 71280 1300
rect 71836 1040 72188 1606
rect 72252 898 72280 1838
rect 73160 1760 73212 1766
rect 73160 1702 73212 1708
rect 73172 1358 73200 1702
rect 73264 1358 73292 2790
rect 74188 2202 74540 3238
rect 74188 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74540 2202
rect 73160 1352 73212 1358
rect 73160 1294 73212 1300
rect 73252 1352 73304 1358
rect 73252 1294 73304 1300
rect 72700 1216 72752 1222
rect 72700 1158 72752 1164
rect 72160 870 72280 898
rect 72160 800 72188 870
rect 72712 800 72740 1158
rect 74188 1114 74540 2150
rect 74188 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74540 1114
rect 74188 1040 74540 1062
rect 64524 734 64736 762
rect 64970 0 65026 800
rect 65522 0 65578 800
rect 66074 0 66130 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68282 0 68338 800
rect 68834 0 68890 800
rect 69386 0 69442 800
rect 69938 0 69994 800
rect 70490 0 70546 800
rect 71042 0 71098 800
rect 71594 0 71650 800
rect 72146 0 72202 800
rect 72698 0 72754 800
<< via2 >>
rect 64216 84532 64272 84588
rect 64296 84532 64352 84588
rect 64376 84532 64432 84588
rect 64456 84532 64512 84588
rect 64216 84452 64272 84508
rect 64296 84452 64352 84508
rect 64376 84452 64432 84508
rect 64456 84452 64512 84508
rect 64216 84372 64272 84428
rect 64296 84372 64352 84428
rect 64376 84372 64432 84428
rect 64456 84372 64512 84428
rect 64216 84292 64272 84348
rect 64296 84292 64352 84348
rect 64376 84292 64432 84348
rect 64456 84292 64512 84348
rect 64216 74532 64272 74588
rect 64296 74532 64352 74588
rect 64376 74532 64432 74588
rect 64456 74532 64512 74588
rect 64216 74452 64272 74508
rect 64296 74452 64352 74508
rect 64376 74452 64432 74508
rect 64456 74452 64512 74508
rect 64216 74372 64272 74428
rect 64296 74372 64352 74428
rect 64376 74372 64432 74428
rect 64456 74372 64512 74428
rect 64216 74292 64272 74348
rect 64296 74292 64352 74348
rect 64376 74292 64432 74348
rect 64456 74292 64512 74348
rect 63498 52572 63500 52592
rect 63500 52572 63552 52592
rect 63552 52572 63554 52592
rect 63498 52536 63554 52572
rect 63498 50260 63500 50280
rect 63500 50260 63552 50280
rect 63552 50260 63554 50280
rect 63498 50224 63554 50260
rect 63406 48769 63408 48784
rect 63408 48769 63460 48784
rect 63460 48769 63462 48784
rect 63406 48728 63462 48769
rect 63498 48061 63500 48104
rect 63500 48061 63552 48104
rect 63552 48061 63554 48104
rect 63498 48048 63554 48061
rect 64216 64532 64272 64588
rect 64296 64532 64352 64588
rect 64376 64532 64432 64588
rect 64456 64532 64512 64588
rect 64216 64452 64272 64508
rect 64296 64452 64352 64508
rect 64376 64452 64432 64508
rect 64456 64452 64512 64508
rect 64216 64372 64272 64428
rect 64296 64372 64352 64428
rect 64376 64372 64432 64428
rect 64456 64372 64512 64428
rect 64216 64292 64272 64348
rect 64296 64292 64352 64348
rect 64376 64292 64432 64348
rect 64456 64292 64512 64348
rect 64216 54532 64272 54588
rect 64296 54532 64352 54588
rect 64376 54532 64432 54588
rect 64456 54532 64512 54588
rect 64216 54452 64272 54508
rect 64296 54452 64352 54508
rect 64376 54452 64432 54508
rect 64456 54452 64512 54508
rect 64216 54372 64272 54428
rect 64296 54372 64352 54428
rect 64376 54372 64432 54428
rect 64456 54372 64512 54428
rect 64216 54292 64272 54348
rect 64296 54292 64352 54348
rect 64376 54292 64432 54348
rect 64456 54292 64512 54348
rect 63866 47676 63868 47696
rect 63868 47676 63920 47696
rect 63920 47676 63922 47696
rect 63866 47640 63922 47676
rect 63682 26152 63738 26208
rect 63498 11736 63554 11792
rect 63406 10648 63462 10704
rect 1864 2180 1920 2236
rect 1944 2180 2000 2236
rect 2024 2180 2080 2236
rect 2104 2180 2160 2236
rect 1864 2100 1920 2156
rect 1944 2100 2000 2156
rect 2024 2100 2080 2156
rect 2104 2100 2160 2156
rect 1864 2020 1920 2076
rect 1944 2020 2000 2076
rect 2024 2020 2080 2076
rect 2104 2020 2160 2076
rect 1864 1940 1920 1996
rect 1944 1940 2000 1996
rect 2024 1940 2080 1996
rect 2104 1940 2160 1996
rect 4216 4532 4272 4588
rect 4296 4532 4352 4588
rect 4376 4532 4432 4588
rect 4456 4532 4512 4588
rect 4216 4452 4272 4508
rect 4296 4452 4352 4508
rect 4376 4452 4432 4508
rect 4456 4452 4512 4508
rect 4216 4378 4272 4428
rect 4296 4378 4352 4428
rect 4376 4378 4432 4428
rect 4456 4378 4512 4428
rect 4216 4372 4262 4378
rect 4262 4372 4272 4378
rect 4296 4372 4326 4378
rect 4326 4372 4338 4378
rect 4338 4372 4352 4378
rect 4376 4372 4390 4378
rect 4390 4372 4402 4378
rect 4402 4372 4432 4378
rect 4456 4372 4466 4378
rect 4466 4372 4512 4378
rect 4216 4326 4262 4348
rect 4262 4326 4272 4348
rect 4296 4326 4326 4348
rect 4326 4326 4338 4348
rect 4338 4326 4352 4348
rect 4376 4326 4390 4348
rect 4390 4326 4402 4348
rect 4402 4326 4432 4348
rect 4456 4326 4466 4348
rect 4466 4326 4512 4348
rect 4216 4292 4272 4326
rect 4296 4292 4352 4326
rect 4376 4292 4432 4326
rect 4456 4292 4512 4326
rect 11864 2180 11920 2236
rect 11944 2180 12000 2236
rect 12024 2180 12080 2236
rect 12104 2180 12160 2236
rect 11864 2100 11920 2156
rect 11944 2100 12000 2156
rect 12024 2100 12080 2156
rect 12104 2100 12160 2156
rect 11864 2020 11920 2076
rect 11944 2020 12000 2076
rect 12024 2020 12080 2076
rect 12104 2020 12160 2076
rect 11864 1940 11920 1996
rect 11944 1940 12000 1996
rect 12024 1940 12080 1996
rect 12104 1940 12160 1996
rect 14216 4532 14272 4588
rect 14296 4532 14352 4588
rect 14376 4532 14432 4588
rect 14456 4532 14512 4588
rect 14216 4452 14272 4508
rect 14296 4452 14352 4508
rect 14376 4452 14432 4508
rect 14456 4452 14512 4508
rect 14216 4378 14272 4428
rect 14296 4378 14352 4428
rect 14376 4378 14432 4428
rect 14456 4378 14512 4428
rect 14216 4372 14262 4378
rect 14262 4372 14272 4378
rect 14296 4372 14326 4378
rect 14326 4372 14338 4378
rect 14338 4372 14352 4378
rect 14376 4372 14390 4378
rect 14390 4372 14402 4378
rect 14402 4372 14432 4378
rect 14456 4372 14466 4378
rect 14466 4372 14512 4378
rect 14216 4326 14262 4348
rect 14262 4326 14272 4348
rect 14296 4326 14326 4348
rect 14326 4326 14338 4348
rect 14338 4326 14352 4348
rect 14376 4326 14390 4348
rect 14390 4326 14402 4348
rect 14402 4326 14432 4348
rect 14456 4326 14466 4348
rect 14466 4326 14512 4348
rect 14216 4292 14272 4326
rect 14296 4292 14352 4326
rect 14376 4292 14432 4326
rect 14456 4292 14512 4326
rect 30286 6840 30342 6896
rect 29642 6704 29698 6760
rect 14738 3304 14794 3360
rect 21864 2180 21920 2236
rect 21944 2180 22000 2236
rect 22024 2180 22080 2236
rect 22104 2180 22160 2236
rect 21864 2100 21920 2156
rect 21944 2100 22000 2156
rect 22024 2100 22080 2156
rect 22104 2100 22160 2156
rect 21864 2020 21920 2076
rect 21944 2020 22000 2076
rect 22024 2020 22080 2076
rect 22104 2020 22160 2076
rect 21864 1940 21920 1996
rect 21944 1940 22000 1996
rect 22024 1940 22080 1996
rect 22104 1940 22160 1996
rect 24216 4532 24272 4588
rect 24296 4532 24352 4588
rect 24376 4532 24432 4588
rect 24456 4532 24512 4588
rect 24216 4452 24272 4508
rect 24296 4452 24352 4508
rect 24376 4452 24432 4508
rect 24456 4452 24512 4508
rect 24216 4378 24272 4428
rect 24296 4378 24352 4428
rect 24376 4378 24432 4428
rect 24456 4378 24512 4428
rect 24216 4372 24262 4378
rect 24262 4372 24272 4378
rect 24296 4372 24326 4378
rect 24326 4372 24338 4378
rect 24338 4372 24352 4378
rect 24376 4372 24390 4378
rect 24390 4372 24402 4378
rect 24402 4372 24432 4378
rect 24456 4372 24466 4378
rect 24466 4372 24512 4378
rect 24216 4326 24262 4348
rect 24262 4326 24272 4348
rect 24296 4326 24326 4348
rect 24326 4326 24338 4348
rect 24338 4326 24352 4348
rect 24376 4326 24390 4348
rect 24390 4326 24402 4348
rect 24402 4326 24432 4348
rect 24456 4326 24466 4348
rect 24466 4326 24512 4348
rect 24216 4292 24272 4326
rect 24296 4292 24352 4326
rect 24376 4292 24432 4326
rect 24456 4292 24512 4326
rect 25870 5888 25926 5944
rect 25870 5108 25872 5128
rect 25872 5108 25924 5128
rect 25924 5108 25926 5128
rect 25870 5072 25926 5108
rect 25502 3476 25504 3496
rect 25504 3476 25556 3496
rect 25556 3476 25558 3496
rect 25502 3440 25558 3476
rect 29274 6568 29330 6624
rect 28446 5344 28502 5400
rect 28170 3440 28226 3496
rect 28998 4936 29054 4992
rect 34058 7520 34114 7576
rect 30838 5228 30894 5264
rect 30838 5208 30840 5228
rect 30840 5208 30892 5228
rect 30892 5208 30894 5228
rect 30378 5108 30380 5128
rect 30380 5108 30432 5128
rect 30432 5108 30434 5128
rect 30378 5072 30434 5108
rect 29642 4936 29698 4992
rect 31298 3984 31354 4040
rect 31298 3440 31354 3496
rect 32218 3032 32274 3088
rect 31864 2180 31920 2236
rect 31944 2180 32000 2236
rect 32024 2180 32080 2236
rect 32104 2180 32160 2236
rect 31864 2100 31920 2156
rect 31944 2100 32000 2156
rect 32024 2100 32080 2156
rect 32104 2100 32160 2156
rect 31864 2020 31920 2076
rect 31944 2020 32000 2076
rect 32024 2020 32080 2076
rect 32104 2020 32160 2076
rect 31864 1940 31920 1996
rect 31944 1940 32000 1996
rect 32024 1940 32080 1996
rect 32104 1940 32160 1996
rect 32770 3596 32826 3632
rect 32770 3576 32772 3596
rect 32772 3576 32824 3596
rect 32824 3576 32826 3596
rect 33230 3440 33286 3496
rect 41050 7656 41106 7712
rect 34216 4532 34272 4588
rect 34296 4532 34352 4588
rect 34376 4532 34432 4588
rect 34456 4532 34512 4588
rect 34216 4452 34272 4508
rect 34296 4452 34352 4508
rect 34376 4452 34432 4508
rect 34456 4452 34512 4508
rect 34216 4378 34272 4428
rect 34296 4378 34352 4428
rect 34376 4378 34432 4428
rect 34456 4378 34512 4428
rect 34216 4372 34262 4378
rect 34262 4372 34272 4378
rect 34296 4372 34326 4378
rect 34326 4372 34338 4378
rect 34338 4372 34352 4378
rect 34376 4372 34390 4378
rect 34390 4372 34402 4378
rect 34402 4372 34432 4378
rect 34456 4372 34466 4378
rect 34466 4372 34512 4378
rect 34216 4326 34262 4348
rect 34262 4326 34272 4348
rect 34296 4326 34326 4348
rect 34326 4326 34338 4348
rect 34338 4326 34352 4348
rect 34376 4326 34390 4348
rect 34390 4326 34402 4348
rect 34402 4326 34432 4348
rect 34456 4326 34466 4348
rect 34466 4326 34512 4348
rect 34216 4292 34272 4326
rect 34296 4292 34352 4326
rect 34376 4292 34432 4326
rect 34456 4292 34512 4326
rect 40406 5752 40462 5808
rect 37002 5636 37058 5672
rect 37002 5616 37004 5636
rect 37004 5616 37056 5636
rect 37056 5616 37058 5636
rect 36082 3596 36138 3632
rect 36082 3576 36084 3596
rect 36084 3576 36136 3596
rect 36136 3576 36138 3596
rect 41694 5616 41750 5672
rect 41864 2180 41920 2236
rect 41944 2180 42000 2236
rect 42024 2180 42080 2236
rect 42104 2180 42160 2236
rect 41864 2100 41920 2156
rect 41944 2100 42000 2156
rect 42024 2100 42080 2156
rect 42104 2100 42160 2156
rect 41864 2020 41920 2076
rect 41944 2020 42000 2076
rect 42024 2020 42080 2076
rect 42104 2020 42160 2076
rect 41864 1940 41920 1996
rect 41944 1940 42000 1996
rect 42024 1940 42080 1996
rect 42104 1940 42160 1996
rect 44638 5888 44694 5944
rect 44086 5108 44088 5128
rect 44088 5108 44140 5128
rect 44140 5108 44142 5128
rect 44086 5072 44142 5108
rect 46018 5480 46074 5536
rect 44216 4532 44272 4588
rect 44296 4532 44352 4588
rect 44376 4532 44432 4588
rect 44456 4532 44512 4588
rect 44216 4452 44272 4508
rect 44296 4452 44352 4508
rect 44376 4452 44432 4508
rect 44456 4452 44512 4508
rect 44216 4378 44272 4428
rect 44296 4378 44352 4428
rect 44376 4378 44432 4428
rect 44456 4378 44512 4428
rect 44216 4372 44262 4378
rect 44262 4372 44272 4378
rect 44296 4372 44326 4378
rect 44326 4372 44338 4378
rect 44338 4372 44352 4378
rect 44376 4372 44390 4378
rect 44390 4372 44402 4378
rect 44402 4372 44432 4378
rect 44456 4372 44466 4378
rect 44466 4372 44512 4378
rect 44216 4326 44262 4348
rect 44262 4326 44272 4348
rect 44296 4326 44326 4348
rect 44326 4326 44338 4348
rect 44338 4326 44352 4348
rect 44376 4326 44390 4348
rect 44390 4326 44402 4348
rect 44402 4326 44432 4348
rect 44456 4326 44466 4348
rect 44466 4326 44512 4348
rect 44216 4292 44272 4326
rect 44296 4292 44352 4326
rect 44376 4292 44432 4326
rect 44456 4292 44512 4326
rect 44730 4936 44786 4992
rect 49514 6024 49570 6080
rect 46662 4800 46718 4856
rect 47582 5072 47638 5128
rect 47858 3304 47914 3360
rect 51864 2180 51920 2236
rect 51944 2180 52000 2236
rect 52024 2180 52080 2236
rect 52104 2180 52160 2236
rect 51864 2100 51920 2156
rect 51944 2100 52000 2156
rect 52024 2100 52080 2156
rect 52104 2100 52160 2156
rect 51864 2020 51920 2076
rect 51944 2020 52000 2076
rect 52024 2020 52080 2076
rect 52104 2020 52160 2076
rect 51864 1940 51920 1996
rect 51944 1940 52000 1996
rect 52024 1940 52080 1996
rect 52104 1940 52160 1996
rect 59558 7792 59614 7848
rect 54216 4532 54272 4588
rect 54296 4532 54352 4588
rect 54376 4532 54432 4588
rect 54456 4532 54512 4588
rect 54216 4452 54272 4508
rect 54296 4452 54352 4508
rect 54376 4452 54432 4508
rect 54456 4452 54512 4508
rect 54216 4378 54272 4428
rect 54296 4378 54352 4428
rect 54376 4378 54432 4428
rect 54456 4378 54512 4428
rect 54216 4372 54262 4378
rect 54262 4372 54272 4378
rect 54296 4372 54326 4378
rect 54326 4372 54338 4378
rect 54338 4372 54352 4378
rect 54376 4372 54390 4378
rect 54390 4372 54402 4378
rect 54402 4372 54432 4378
rect 54456 4372 54466 4378
rect 54466 4372 54512 4378
rect 54216 4326 54262 4348
rect 54262 4326 54272 4348
rect 54296 4326 54326 4348
rect 54326 4326 54338 4348
rect 54338 4326 54352 4348
rect 54376 4326 54390 4348
rect 54390 4326 54402 4348
rect 54402 4326 54432 4348
rect 54456 4326 54466 4348
rect 54466 4326 54512 4348
rect 54216 4292 54272 4326
rect 54296 4292 54352 4326
rect 54376 4292 54432 4326
rect 54456 4292 54512 4326
rect 59174 7384 59230 7440
rect 56506 6296 56562 6352
rect 55770 6160 55826 6216
rect 55770 5752 55826 5808
rect 57518 6024 57574 6080
rect 58162 6024 58218 6080
rect 55862 5480 55918 5536
rect 55862 5072 55918 5128
rect 59634 6976 59690 7032
rect 60922 5480 60978 5536
rect 61014 4120 61070 4176
rect 61474 4120 61530 4176
rect 63498 7248 63554 7304
rect 62762 6024 62818 6080
rect 63130 6024 63186 6080
rect 62946 5752 63002 5808
rect 63406 5752 63462 5808
rect 63130 5344 63186 5400
rect 63406 5344 63462 5400
rect 63774 16496 63830 16552
rect 63590 6296 63646 6352
rect 63406 4800 63462 4856
rect 63590 4800 63646 4856
rect 61864 2180 61920 2236
rect 61944 2180 62000 2236
rect 62024 2180 62080 2236
rect 62104 2180 62160 2236
rect 61864 2100 61920 2156
rect 61944 2100 62000 2156
rect 62024 2100 62080 2156
rect 62104 2100 62160 2156
rect 61864 2020 61920 2076
rect 61944 2020 62000 2076
rect 62024 2020 62080 2076
rect 62104 2020 62160 2076
rect 61864 1940 61920 1996
rect 61944 1940 62000 1996
rect 62024 1940 62080 1996
rect 62104 1940 62160 1996
rect 64216 44532 64272 44588
rect 64296 44532 64352 44588
rect 64376 44532 64432 44588
rect 64456 44532 64512 44588
rect 64216 44452 64272 44508
rect 64296 44452 64352 44508
rect 64376 44452 64432 44508
rect 64456 44452 64512 44508
rect 64216 44372 64272 44428
rect 64296 44372 64352 44428
rect 64376 44372 64432 44428
rect 64456 44372 64512 44428
rect 64216 44292 64272 44348
rect 64296 44292 64352 44348
rect 64376 44292 64432 44348
rect 64456 44292 64512 44348
rect 64216 34532 64272 34588
rect 64296 34532 64352 34588
rect 64376 34532 64432 34588
rect 64456 34532 64512 34588
rect 64216 34452 64272 34508
rect 64296 34452 64352 34508
rect 64376 34452 64432 34508
rect 64456 34452 64512 34508
rect 64216 34372 64272 34428
rect 64296 34372 64352 34428
rect 64376 34372 64432 34428
rect 64456 34372 64512 34428
rect 64216 34292 64272 34348
rect 64296 34292 64352 34348
rect 64376 34292 64432 34348
rect 64456 34292 64512 34348
rect 64216 24532 64272 24588
rect 64296 24532 64352 24588
rect 64376 24532 64432 24588
rect 64456 24532 64512 24588
rect 64216 24452 64272 24508
rect 64296 24452 64352 24508
rect 64376 24452 64432 24508
rect 64456 24452 64512 24508
rect 64216 24372 64272 24428
rect 64296 24372 64352 24428
rect 64376 24372 64432 24428
rect 64456 24372 64512 24428
rect 64216 24292 64272 24348
rect 64296 24292 64352 24348
rect 64376 24292 64432 24348
rect 64456 24292 64512 24348
rect 64216 14532 64272 14588
rect 64296 14532 64352 14588
rect 64376 14532 64432 14588
rect 64456 14532 64512 14588
rect 64216 14452 64272 14508
rect 64296 14452 64352 14508
rect 64376 14452 64432 14508
rect 64456 14452 64512 14508
rect 64216 14372 64272 14428
rect 64296 14372 64352 14428
rect 64376 14372 64432 14428
rect 64456 14372 64512 14428
rect 64216 14292 64272 14348
rect 64296 14292 64352 14348
rect 64376 14292 64432 14348
rect 64456 14292 64512 14348
rect 64050 11192 64106 11248
rect 64050 7928 64106 7984
rect 64216 4532 64272 4588
rect 64296 4532 64352 4588
rect 64376 4532 64432 4588
rect 64456 4532 64512 4588
rect 64216 4452 64272 4508
rect 64296 4452 64352 4508
rect 64376 4452 64432 4508
rect 64456 4452 64512 4508
rect 64216 4378 64272 4428
rect 64296 4378 64352 4428
rect 64376 4378 64432 4428
rect 64456 4378 64512 4428
rect 64216 4372 64262 4378
rect 64262 4372 64272 4378
rect 64296 4372 64326 4378
rect 64326 4372 64338 4378
rect 64338 4372 64352 4378
rect 64376 4372 64390 4378
rect 64390 4372 64402 4378
rect 64402 4372 64432 4378
rect 64456 4372 64466 4378
rect 64466 4372 64512 4378
rect 64216 4326 64262 4348
rect 64262 4326 64272 4348
rect 64296 4326 64326 4348
rect 64326 4326 64338 4348
rect 64338 4326 64352 4348
rect 64376 4326 64390 4348
rect 64390 4326 64402 4348
rect 64402 4326 64432 4348
rect 64456 4326 64466 4348
rect 64466 4326 64512 4348
rect 64216 4292 64272 4326
rect 64296 4292 64352 4326
rect 64376 4292 64432 4326
rect 64456 4292 64512 4326
rect 64970 40840 65026 40896
rect 64970 38836 64972 38856
rect 64972 38836 65024 38856
rect 65024 38836 65026 38856
rect 64970 38800 65026 38836
rect 65522 34720 65578 34776
rect 65614 33224 65670 33280
rect 64878 12724 64880 12744
rect 64880 12724 64932 12744
rect 64932 12724 64934 12744
rect 64878 12688 64934 12724
rect 64878 12552 64934 12608
rect 64878 11736 64934 11792
rect 64878 6296 64934 6352
rect 64786 5888 64842 5944
rect 64970 5480 65026 5536
rect 64878 3032 64934 3088
rect 66074 6432 66130 6488
rect 66442 23432 66498 23488
rect 66442 22344 66498 22400
rect 67178 7384 67234 7440
rect 67362 26424 67418 26480
rect 67546 26016 67602 26072
rect 67638 23604 67640 23624
rect 67640 23604 67692 23624
rect 67692 23604 67694 23624
rect 67638 23568 67694 23604
rect 69018 5752 69074 5808
rect 69110 5344 69166 5400
rect 71864 82180 71920 82236
rect 71944 82180 72000 82236
rect 72024 82180 72080 82236
rect 72104 82180 72160 82236
rect 71864 82118 71910 82156
rect 71910 82118 71920 82156
rect 71944 82118 71974 82156
rect 71974 82118 71986 82156
rect 71986 82118 72000 82156
rect 72024 82118 72038 82156
rect 72038 82118 72050 82156
rect 72050 82118 72080 82156
rect 72104 82118 72114 82156
rect 72114 82118 72160 82156
rect 71864 82100 71920 82118
rect 71944 82100 72000 82118
rect 72024 82100 72080 82118
rect 72104 82100 72160 82118
rect 71864 82020 71920 82076
rect 71944 82020 72000 82076
rect 72024 82020 72080 82076
rect 72104 82020 72160 82076
rect 71864 81940 71920 81996
rect 71944 81940 72000 81996
rect 72024 81940 72080 81996
rect 72104 81940 72160 81996
rect 71864 72180 71920 72236
rect 71944 72180 72000 72236
rect 72024 72180 72080 72236
rect 72104 72180 72160 72236
rect 71864 72100 71920 72156
rect 71944 72100 72000 72156
rect 72024 72100 72080 72156
rect 72104 72100 72160 72156
rect 71864 72020 71920 72076
rect 71944 72020 72000 72076
rect 72024 72020 72080 72076
rect 72104 72020 72160 72076
rect 71864 71940 71920 71996
rect 71944 71940 72000 71996
rect 72024 71940 72080 71996
rect 72104 71940 72160 71996
rect 71864 62180 71920 62236
rect 71944 62180 72000 62236
rect 72024 62180 72080 62236
rect 72104 62180 72160 62236
rect 71864 62100 71920 62156
rect 71944 62100 72000 62156
rect 72024 62100 72080 62156
rect 72104 62100 72160 62156
rect 71864 62020 71920 62076
rect 71944 62020 72000 62076
rect 72024 62020 72080 62076
rect 72104 62020 72160 62076
rect 71864 61940 71920 61996
rect 71944 61940 72000 61996
rect 72024 61940 72080 61996
rect 72104 61940 72160 61996
rect 70490 5208 70546 5264
rect 71864 52180 71920 52236
rect 71944 52180 72000 52236
rect 72024 52180 72080 52236
rect 72104 52180 72160 52236
rect 71864 52100 71920 52156
rect 71944 52100 72000 52156
rect 72024 52100 72080 52156
rect 72104 52100 72160 52156
rect 71864 52020 71920 52076
rect 71944 52020 72000 52076
rect 72024 52020 72080 52076
rect 72104 52020 72160 52076
rect 71864 51940 71920 51996
rect 71944 51940 72000 51996
rect 72024 51940 72080 51996
rect 72104 51940 72160 51996
rect 71864 42180 71920 42236
rect 71944 42180 72000 42236
rect 72024 42180 72080 42236
rect 72104 42180 72160 42236
rect 71864 42100 71920 42156
rect 71944 42100 72000 42156
rect 72024 42100 72080 42156
rect 72104 42100 72160 42156
rect 71864 42020 71920 42076
rect 71944 42020 72000 42076
rect 72024 42020 72080 42076
rect 72104 42020 72160 42076
rect 71864 41940 71920 41996
rect 71944 41940 72000 41996
rect 72024 41940 72080 41996
rect 72104 41940 72160 41996
rect 71864 32180 71920 32236
rect 71944 32180 72000 32236
rect 72024 32180 72080 32236
rect 72104 32180 72160 32236
rect 71864 32122 71920 32156
rect 71944 32122 72000 32156
rect 72024 32122 72080 32156
rect 72104 32122 72160 32156
rect 71864 32100 71910 32122
rect 71910 32100 71920 32122
rect 71944 32100 71974 32122
rect 71974 32100 71986 32122
rect 71986 32100 72000 32122
rect 72024 32100 72038 32122
rect 72038 32100 72050 32122
rect 72050 32100 72080 32122
rect 72104 32100 72114 32122
rect 72114 32100 72160 32122
rect 71864 32070 71910 32076
rect 71910 32070 71920 32076
rect 71944 32070 71974 32076
rect 71974 32070 71986 32076
rect 71986 32070 72000 32076
rect 72024 32070 72038 32076
rect 72038 32070 72050 32076
rect 72050 32070 72080 32076
rect 72104 32070 72114 32076
rect 72114 32070 72160 32076
rect 71864 32020 71920 32070
rect 71944 32020 72000 32070
rect 72024 32020 72080 32070
rect 72104 32020 72160 32070
rect 71864 31940 71920 31996
rect 71944 31940 72000 31996
rect 72024 31940 72080 31996
rect 72104 31940 72160 31996
rect 71864 22180 71920 22236
rect 71944 22180 72000 22236
rect 72024 22180 72080 22236
rect 72104 22180 72160 22236
rect 71864 22100 71920 22156
rect 71944 22100 72000 22156
rect 72024 22100 72080 22156
rect 72104 22100 72160 22156
rect 71864 22020 71920 22076
rect 71944 22020 72000 22076
rect 72024 22020 72080 22076
rect 72104 22020 72160 22076
rect 71864 21940 71920 21996
rect 71944 21940 72000 21996
rect 72024 21940 72080 21996
rect 72104 21940 72160 21996
rect 71864 12180 71920 12236
rect 71944 12180 72000 12236
rect 72024 12180 72080 12236
rect 72104 12180 72160 12236
rect 71864 12100 71920 12156
rect 71944 12100 72000 12156
rect 72024 12100 72080 12156
rect 72104 12100 72160 12156
rect 71864 12020 71920 12076
rect 71944 12020 72000 12076
rect 72024 12020 72080 12076
rect 72104 12020 72160 12076
rect 71864 11940 71920 11996
rect 71944 11940 72000 11996
rect 72024 11940 72080 11996
rect 72104 11940 72160 11996
rect 74216 84532 74272 84588
rect 74296 84532 74352 84588
rect 74376 84532 74432 84588
rect 74456 84532 74512 84588
rect 74216 84452 74272 84508
rect 74296 84452 74352 84508
rect 74376 84452 74432 84508
rect 74456 84452 74512 84508
rect 74216 84372 74272 84428
rect 74296 84372 74352 84428
rect 74376 84372 74432 84428
rect 74456 84372 74512 84428
rect 74216 84292 74272 84348
rect 74296 84292 74352 84348
rect 74376 84292 74432 84348
rect 74456 84292 74512 84348
rect 74216 74532 74272 74588
rect 74296 74532 74352 74588
rect 74376 74532 74432 74588
rect 74456 74532 74512 74588
rect 74216 74452 74272 74508
rect 74296 74452 74352 74508
rect 74376 74452 74432 74508
rect 74456 74452 74512 74508
rect 74216 74372 74272 74428
rect 74296 74372 74352 74428
rect 74376 74372 74432 74428
rect 74456 74372 74512 74428
rect 74216 74292 74272 74348
rect 74296 74292 74352 74348
rect 74376 74292 74432 74348
rect 74456 74292 74512 74348
rect 74216 64532 74272 64588
rect 74296 64532 74352 64588
rect 74376 64532 74432 64588
rect 74456 64532 74512 64588
rect 74216 64452 74272 64508
rect 74296 64452 74352 64508
rect 74376 64452 74432 64508
rect 74456 64452 74512 64508
rect 74216 64372 74272 64428
rect 74296 64372 74352 64428
rect 74376 64372 74432 64428
rect 74456 64372 74512 64428
rect 74216 64292 74272 64348
rect 74296 64292 74352 64348
rect 74376 64292 74432 64348
rect 74456 64292 74512 64348
rect 74216 54532 74272 54588
rect 74296 54532 74352 54588
rect 74376 54532 74432 54588
rect 74456 54532 74512 54588
rect 74216 54452 74272 54508
rect 74296 54452 74352 54508
rect 74376 54452 74432 54508
rect 74456 54452 74512 54508
rect 74216 54426 74272 54428
rect 74296 54426 74352 54428
rect 74376 54426 74432 54428
rect 74456 54426 74512 54428
rect 74216 54374 74262 54426
rect 74262 54374 74272 54426
rect 74296 54374 74326 54426
rect 74326 54374 74338 54426
rect 74338 54374 74352 54426
rect 74376 54374 74390 54426
rect 74390 54374 74402 54426
rect 74402 54374 74432 54426
rect 74456 54374 74466 54426
rect 74466 54374 74512 54426
rect 74216 54372 74272 54374
rect 74296 54372 74352 54374
rect 74376 54372 74432 54374
rect 74456 54372 74512 54374
rect 74216 54292 74272 54348
rect 74296 54292 74352 54348
rect 74376 54292 74432 54348
rect 74456 54292 74512 54348
rect 74216 44582 74262 44588
rect 74262 44582 74272 44588
rect 74296 44582 74326 44588
rect 74326 44582 74338 44588
rect 74338 44582 74352 44588
rect 74376 44582 74390 44588
rect 74390 44582 74402 44588
rect 74402 44582 74432 44588
rect 74456 44582 74466 44588
rect 74466 44582 74512 44588
rect 74216 44532 74272 44582
rect 74296 44532 74352 44582
rect 74376 44532 74432 44582
rect 74456 44532 74512 44582
rect 74216 44452 74272 44508
rect 74296 44452 74352 44508
rect 74376 44452 74432 44508
rect 74456 44452 74512 44508
rect 74216 44372 74272 44428
rect 74296 44372 74352 44428
rect 74376 44372 74432 44428
rect 74456 44372 74512 44428
rect 74216 44292 74272 44348
rect 74296 44292 74352 44348
rect 74376 44292 74432 44348
rect 74456 44292 74512 44348
rect 74216 34532 74272 34588
rect 74296 34532 74352 34588
rect 74376 34532 74432 34588
rect 74456 34532 74512 34588
rect 74216 34452 74272 34508
rect 74296 34452 74352 34508
rect 74376 34452 74432 34508
rect 74456 34452 74512 34508
rect 74216 34372 74272 34428
rect 74296 34372 74352 34428
rect 74376 34372 74432 34428
rect 74456 34372 74512 34428
rect 74216 34292 74272 34348
rect 74296 34292 74352 34348
rect 74376 34292 74432 34348
rect 74456 34292 74512 34348
rect 74216 24532 74272 24588
rect 74296 24532 74352 24588
rect 74376 24532 74432 24588
rect 74456 24532 74512 24588
rect 74216 24452 74272 24508
rect 74296 24452 74352 24508
rect 74376 24452 74432 24508
rect 74456 24452 74512 24508
rect 74216 24372 74272 24428
rect 74296 24372 74352 24428
rect 74376 24372 74432 24428
rect 74456 24372 74512 24428
rect 74216 24292 74272 24348
rect 74296 24292 74352 24348
rect 74376 24292 74432 24348
rect 74456 24292 74512 24348
rect 74216 14532 74272 14588
rect 74296 14532 74352 14588
rect 74376 14532 74432 14588
rect 74456 14532 74512 14588
rect 74216 14452 74272 14508
rect 74296 14452 74352 14508
rect 74376 14452 74432 14508
rect 74456 14452 74512 14508
rect 74216 14372 74272 14428
rect 74296 14372 74352 14428
rect 74376 14372 74432 14428
rect 74456 14372 74512 14428
rect 74216 14292 74272 14348
rect 74296 14292 74352 14348
rect 74376 14292 74432 14348
rect 74456 14292 74512 14348
rect 74216 4532 74272 4588
rect 74296 4532 74352 4588
rect 74376 4532 74432 4588
rect 74456 4532 74512 4588
rect 74216 4452 74272 4508
rect 74296 4452 74352 4508
rect 74376 4452 74432 4508
rect 74456 4452 74512 4508
rect 74216 4378 74272 4428
rect 74296 4378 74352 4428
rect 74376 4378 74432 4428
rect 74456 4378 74512 4428
rect 74216 4372 74262 4378
rect 74262 4372 74272 4378
rect 74296 4372 74326 4378
rect 74326 4372 74338 4378
rect 74338 4372 74352 4378
rect 74376 4372 74390 4378
rect 74390 4372 74402 4378
rect 74402 4372 74432 4378
rect 74456 4372 74466 4378
rect 74466 4372 74512 4378
rect 74216 4326 74262 4348
rect 74262 4326 74272 4348
rect 74296 4326 74326 4348
rect 74326 4326 74338 4348
rect 74338 4326 74352 4348
rect 74376 4326 74390 4348
rect 74390 4326 74402 4348
rect 74402 4326 74432 4348
rect 74456 4326 74466 4348
rect 74466 4326 74512 4348
rect 74216 4292 74272 4326
rect 74296 4292 74352 4326
rect 74376 4292 74432 4326
rect 74456 4292 74512 4326
rect 71864 2180 71920 2236
rect 71944 2180 72000 2236
rect 72024 2180 72080 2236
rect 72104 2180 72160 2236
rect 71864 2100 71920 2156
rect 71944 2100 72000 2156
rect 72024 2100 72080 2156
rect 72104 2100 72160 2156
rect 71864 2020 71920 2076
rect 71944 2020 72000 2076
rect 72024 2020 72080 2076
rect 72104 2020 72160 2076
rect 71864 1940 71920 1996
rect 71944 1940 72000 1996
rect 72024 1940 72080 1996
rect 72104 1940 72160 1996
<< metal3 >>
rect 964 84592 75028 84616
rect 964 84528 4740 84592
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84528 10740 84592
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84528 16740 84592
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84528 17140 84592
rect 17204 84528 17220 84592
rect 17284 84528 22740 84592
rect 22804 84528 22820 84592
rect 22884 84528 22900 84592
rect 22964 84528 22980 84592
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84528 28740 84592
rect 28804 84528 28820 84592
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84528 34740 84592
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84528 40740 84592
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84528 46740 84592
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84528 52740 84592
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84528 58740 84592
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84528 59060 84592
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84588 64740 84592
rect 59284 84532 64216 84588
rect 64272 84532 64296 84588
rect 64352 84532 64376 84588
rect 64432 84532 64456 84588
rect 64512 84532 64740 84588
rect 59284 84528 64740 84532
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84588 75028 84592
rect 71284 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 75028 84588
rect 71284 84528 75028 84532
rect 964 84512 75028 84528
rect 964 84448 4740 84512
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84448 10740 84512
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84448 16740 84512
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84448 17140 84512
rect 17204 84448 17220 84512
rect 17284 84448 22740 84512
rect 22804 84448 22820 84512
rect 22884 84448 22900 84512
rect 22964 84448 22980 84512
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84448 28740 84512
rect 28804 84448 28820 84512
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84448 34740 84512
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84448 40740 84512
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84448 46740 84512
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84448 52740 84512
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84448 58740 84512
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84448 59060 84512
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84508 64740 84512
rect 59284 84452 64216 84508
rect 64272 84452 64296 84508
rect 64352 84452 64376 84508
rect 64432 84452 64456 84508
rect 64512 84452 64740 84508
rect 59284 84448 64740 84452
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84508 75028 84512
rect 71284 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 75028 84508
rect 71284 84448 75028 84452
rect 964 84432 75028 84448
rect 964 84368 4740 84432
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84368 10740 84432
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84368 16740 84432
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84368 17140 84432
rect 17204 84368 17220 84432
rect 17284 84368 22740 84432
rect 22804 84368 22820 84432
rect 22884 84368 22900 84432
rect 22964 84368 22980 84432
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84368 28740 84432
rect 28804 84368 28820 84432
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84368 34740 84432
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84368 40740 84432
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84368 46740 84432
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84368 52740 84432
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84368 58740 84432
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84368 59060 84432
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84428 64740 84432
rect 59284 84372 64216 84428
rect 64272 84372 64296 84428
rect 64352 84372 64376 84428
rect 64432 84372 64456 84428
rect 64512 84372 64740 84428
rect 59284 84368 64740 84372
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84428 75028 84432
rect 71284 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 75028 84428
rect 71284 84368 75028 84372
rect 964 84352 75028 84368
rect 964 84288 4740 84352
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84288 10740 84352
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84288 16740 84352
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84288 17140 84352
rect 17204 84288 17220 84352
rect 17284 84288 22740 84352
rect 22804 84288 22820 84352
rect 22884 84288 22900 84352
rect 22964 84288 22980 84352
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84288 28740 84352
rect 28804 84288 28820 84352
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84288 34740 84352
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84288 40740 84352
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84288 46740 84352
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84288 52740 84352
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84288 58740 84352
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84288 59060 84352
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84348 64740 84352
rect 59284 84292 64216 84348
rect 64272 84292 64296 84348
rect 64352 84292 64376 84348
rect 64432 84292 64456 84348
rect 64512 84292 64740 84348
rect 59284 84288 64740 84292
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84348 75028 84352
rect 71284 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 75028 84348
rect 71284 84288 75028 84292
rect 964 84264 75028 84288
rect 964 82240 75028 82264
rect 964 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82176 2220 82240
rect 2284 82176 7740 82240
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82176 13740 82240
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82176 14220 82240
rect 14284 82176 19740 82240
rect 19804 82176 19820 82240
rect 19884 82176 19900 82240
rect 19964 82176 19980 82240
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82176 25740 82240
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82176 31740 82240
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82176 37740 82240
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82176 43740 82240
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82176 49740 82240
rect 49804 82176 49820 82240
rect 49884 82176 49900 82240
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82176 55740 82240
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82176 61740 82240
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82176 67740 82240
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82236 73740 82240
rect 68284 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 73740 82236
rect 68284 82176 73740 82180
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 75028 82240
rect 964 82160 75028 82176
rect 964 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82096 2220 82160
rect 2284 82096 7740 82160
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82096 13740 82160
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82096 14220 82160
rect 14284 82096 19740 82160
rect 19804 82096 19820 82160
rect 19884 82096 19900 82160
rect 19964 82096 19980 82160
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82096 25740 82160
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82096 31740 82160
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82096 37740 82160
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82096 43740 82160
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82096 49740 82160
rect 49804 82096 49820 82160
rect 49884 82096 49900 82160
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82096 55740 82160
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82096 61740 82160
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82096 67740 82160
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82156 73740 82160
rect 68284 82100 71864 82156
rect 71920 82100 71944 82156
rect 72000 82100 72024 82156
rect 72080 82100 72104 82156
rect 72160 82100 73740 82156
rect 68284 82096 73740 82100
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 75028 82160
rect 964 82080 75028 82096
rect 964 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82016 2220 82080
rect 2284 82016 7740 82080
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82016 13740 82080
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82016 14220 82080
rect 14284 82016 19740 82080
rect 19804 82016 19820 82080
rect 19884 82016 19900 82080
rect 19964 82016 19980 82080
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82016 25740 82080
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82016 31740 82080
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82016 37740 82080
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82016 43740 82080
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82016 49740 82080
rect 49804 82016 49820 82080
rect 49884 82016 49900 82080
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82016 55740 82080
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82016 61740 82080
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82016 67740 82080
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82076 73740 82080
rect 68284 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 73740 82076
rect 68284 82016 73740 82020
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 75028 82080
rect 964 82000 75028 82016
rect 964 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81936 2220 82000
rect 2284 81936 7740 82000
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81936 13740 82000
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81936 14220 82000
rect 14284 81936 19740 82000
rect 19804 81936 19820 82000
rect 19884 81936 19900 82000
rect 19964 81936 19980 82000
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81936 25740 82000
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81936 31740 82000
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81936 37740 82000
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81936 43740 82000
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81936 49740 82000
rect 49804 81936 49820 82000
rect 49884 81936 49900 82000
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81936 55740 82000
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81936 61740 82000
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81936 67740 82000
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81996 73740 82000
rect 68284 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 73740 81996
rect 68284 81936 73740 81940
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 75028 82000
rect 964 81912 75028 81936
rect 964 74592 75028 74616
rect 964 74528 4740 74592
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74528 10740 74592
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74528 16740 74592
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74528 17140 74592
rect 17204 74528 17220 74592
rect 17284 74528 22740 74592
rect 22804 74528 22820 74592
rect 22884 74528 22900 74592
rect 22964 74528 22980 74592
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74528 28740 74592
rect 28804 74528 28820 74592
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74528 34740 74592
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74528 40740 74592
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74528 46740 74592
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74528 52740 74592
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74528 58740 74592
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74528 59060 74592
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74588 64740 74592
rect 59284 74532 64216 74588
rect 64272 74532 64296 74588
rect 64352 74532 64376 74588
rect 64432 74532 64456 74588
rect 64512 74532 64740 74588
rect 59284 74528 64740 74532
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74588 75028 74592
rect 71284 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 75028 74588
rect 71284 74528 75028 74532
rect 964 74512 75028 74528
rect 964 74448 4740 74512
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74448 10740 74512
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74448 16740 74512
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74448 17140 74512
rect 17204 74448 17220 74512
rect 17284 74448 22740 74512
rect 22804 74448 22820 74512
rect 22884 74448 22900 74512
rect 22964 74448 22980 74512
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74448 28740 74512
rect 28804 74448 28820 74512
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74448 34740 74512
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74448 40740 74512
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74448 46740 74512
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74448 52740 74512
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74448 58740 74512
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74448 59060 74512
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74508 64740 74512
rect 59284 74452 64216 74508
rect 64272 74452 64296 74508
rect 64352 74452 64376 74508
rect 64432 74452 64456 74508
rect 64512 74452 64740 74508
rect 59284 74448 64740 74452
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74508 75028 74512
rect 71284 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 75028 74508
rect 71284 74448 75028 74452
rect 964 74432 75028 74448
rect 964 74368 4740 74432
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74368 10740 74432
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74368 16740 74432
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74368 17140 74432
rect 17204 74368 17220 74432
rect 17284 74368 22740 74432
rect 22804 74368 22820 74432
rect 22884 74368 22900 74432
rect 22964 74368 22980 74432
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74368 28740 74432
rect 28804 74368 28820 74432
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74368 34740 74432
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74368 40740 74432
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74368 46740 74432
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74368 52740 74432
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74368 58740 74432
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74368 59060 74432
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74428 64740 74432
rect 59284 74372 64216 74428
rect 64272 74372 64296 74428
rect 64352 74372 64376 74428
rect 64432 74372 64456 74428
rect 64512 74372 64740 74428
rect 59284 74368 64740 74372
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74428 75028 74432
rect 71284 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 75028 74428
rect 71284 74368 75028 74372
rect 964 74352 75028 74368
rect 964 74288 4740 74352
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74288 10740 74352
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74288 16740 74352
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74288 17140 74352
rect 17204 74288 17220 74352
rect 17284 74288 22740 74352
rect 22804 74288 22820 74352
rect 22884 74288 22900 74352
rect 22964 74288 22980 74352
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74288 28740 74352
rect 28804 74288 28820 74352
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74288 34740 74352
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74288 40740 74352
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74288 46740 74352
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74288 52740 74352
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74288 58740 74352
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74288 59060 74352
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74348 64740 74352
rect 59284 74292 64216 74348
rect 64272 74292 64296 74348
rect 64352 74292 64376 74348
rect 64432 74292 64456 74348
rect 64512 74292 64740 74348
rect 59284 74288 64740 74292
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74348 75028 74352
rect 71284 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 75028 74348
rect 71284 74288 75028 74292
rect 964 74264 75028 74288
rect 964 72240 75028 72264
rect 964 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72176 2220 72240
rect 2284 72176 7740 72240
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72176 13740 72240
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72176 14220 72240
rect 14284 72176 19740 72240
rect 19804 72176 19820 72240
rect 19884 72176 19900 72240
rect 19964 72176 19980 72240
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72176 25740 72240
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72176 31740 72240
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72176 37740 72240
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72176 43740 72240
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72176 49740 72240
rect 49804 72176 49820 72240
rect 49884 72176 49900 72240
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72176 55740 72240
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72176 61740 72240
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72176 67740 72240
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72236 73740 72240
rect 68284 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 73740 72236
rect 68284 72176 73740 72180
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 75028 72240
rect 964 72160 75028 72176
rect 964 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72096 2220 72160
rect 2284 72096 7740 72160
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72096 13740 72160
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72096 14220 72160
rect 14284 72096 19740 72160
rect 19804 72096 19820 72160
rect 19884 72096 19900 72160
rect 19964 72096 19980 72160
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72096 25740 72160
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72096 31740 72160
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72096 37740 72160
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72096 43740 72160
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72096 49740 72160
rect 49804 72096 49820 72160
rect 49884 72096 49900 72160
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72096 55740 72160
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72096 61740 72160
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72096 67740 72160
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72156 73740 72160
rect 68284 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 73740 72156
rect 68284 72096 73740 72100
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 75028 72160
rect 964 72080 75028 72096
rect 964 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72016 2220 72080
rect 2284 72016 7740 72080
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72016 13740 72080
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72016 14220 72080
rect 14284 72016 19740 72080
rect 19804 72016 19820 72080
rect 19884 72016 19900 72080
rect 19964 72016 19980 72080
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72016 25740 72080
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72016 31740 72080
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72016 37740 72080
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72016 43740 72080
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72016 49740 72080
rect 49804 72016 49820 72080
rect 49884 72016 49900 72080
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72016 55740 72080
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72016 61740 72080
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72016 67740 72080
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72076 73740 72080
rect 68284 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 73740 72076
rect 68284 72016 73740 72020
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 75028 72080
rect 964 72000 75028 72016
rect 964 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71936 2220 72000
rect 2284 71936 7740 72000
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71936 13740 72000
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71936 14220 72000
rect 14284 71936 19740 72000
rect 19804 71936 19820 72000
rect 19884 71936 19900 72000
rect 19964 71936 19980 72000
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71936 25740 72000
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71936 31740 72000
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71936 37740 72000
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71936 43740 72000
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71936 49740 72000
rect 49804 71936 49820 72000
rect 49884 71936 49900 72000
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71936 55740 72000
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71936 61740 72000
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71936 67740 72000
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71996 73740 72000
rect 68284 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 73740 71996
rect 68284 71936 73740 71940
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 75028 72000
rect 964 71912 75028 71936
rect 964 64592 75028 64616
rect 964 64528 4740 64592
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64528 10740 64592
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64528 16740 64592
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64528 17140 64592
rect 17204 64528 17220 64592
rect 17284 64528 22740 64592
rect 22804 64528 22820 64592
rect 22884 64528 22900 64592
rect 22964 64528 22980 64592
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64528 28740 64592
rect 28804 64528 28820 64592
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64528 34740 64592
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64528 40740 64592
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64528 46740 64592
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64528 52740 64592
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64528 58740 64592
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64528 59060 64592
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64588 64740 64592
rect 59284 64532 64216 64588
rect 64272 64532 64296 64588
rect 64352 64532 64376 64588
rect 64432 64532 64456 64588
rect 64512 64532 64740 64588
rect 59284 64528 64740 64532
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64588 75028 64592
rect 71284 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 75028 64588
rect 71284 64528 75028 64532
rect 964 64512 75028 64528
rect 964 64448 4740 64512
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64448 10740 64512
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64448 16740 64512
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64448 17140 64512
rect 17204 64448 17220 64512
rect 17284 64448 22740 64512
rect 22804 64448 22820 64512
rect 22884 64448 22900 64512
rect 22964 64448 22980 64512
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64448 28740 64512
rect 28804 64448 28820 64512
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64448 34740 64512
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64448 40740 64512
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64448 46740 64512
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64448 52740 64512
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64448 58740 64512
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64448 59060 64512
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64508 64740 64512
rect 59284 64452 64216 64508
rect 64272 64452 64296 64508
rect 64352 64452 64376 64508
rect 64432 64452 64456 64508
rect 64512 64452 64740 64508
rect 59284 64448 64740 64452
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64508 75028 64512
rect 71284 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 75028 64508
rect 71284 64448 75028 64452
rect 964 64432 75028 64448
rect 964 64368 4740 64432
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64368 10740 64432
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64368 16740 64432
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64368 17140 64432
rect 17204 64368 17220 64432
rect 17284 64368 22740 64432
rect 22804 64368 22820 64432
rect 22884 64368 22900 64432
rect 22964 64368 22980 64432
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64368 28740 64432
rect 28804 64368 28820 64432
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64368 34740 64432
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64368 40740 64432
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64368 46740 64432
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64368 52740 64432
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64368 58740 64432
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64368 59060 64432
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64428 64740 64432
rect 59284 64372 64216 64428
rect 64272 64372 64296 64428
rect 64352 64372 64376 64428
rect 64432 64372 64456 64428
rect 64512 64372 64740 64428
rect 59284 64368 64740 64372
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64428 75028 64432
rect 71284 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 75028 64428
rect 71284 64368 75028 64372
rect 964 64352 75028 64368
rect 964 64288 4740 64352
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64288 10740 64352
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64288 16740 64352
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64288 17140 64352
rect 17204 64288 17220 64352
rect 17284 64288 22740 64352
rect 22804 64288 22820 64352
rect 22884 64288 22900 64352
rect 22964 64288 22980 64352
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64288 28740 64352
rect 28804 64288 28820 64352
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64288 34740 64352
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64288 40740 64352
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64288 46740 64352
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64288 52740 64352
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64288 58740 64352
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64288 59060 64352
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64348 64740 64352
rect 59284 64292 64216 64348
rect 64272 64292 64296 64348
rect 64352 64292 64376 64348
rect 64432 64292 64456 64348
rect 64512 64292 64740 64348
rect 59284 64288 64740 64292
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64348 75028 64352
rect 71284 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 75028 64348
rect 71284 64288 75028 64292
rect 964 64264 75028 64288
rect 964 62240 75028 62264
rect 964 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62176 2220 62240
rect 2284 62176 7740 62240
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62176 13740 62240
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62176 14220 62240
rect 14284 62176 19740 62240
rect 19804 62176 19820 62240
rect 19884 62176 19900 62240
rect 19964 62176 19980 62240
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62176 25740 62240
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62176 31740 62240
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62176 37740 62240
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62176 43740 62240
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62176 49740 62240
rect 49804 62176 49820 62240
rect 49884 62176 49900 62240
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62176 55740 62240
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62176 61740 62240
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62176 67740 62240
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62236 73740 62240
rect 68284 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 73740 62236
rect 68284 62176 73740 62180
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 75028 62240
rect 964 62160 75028 62176
rect 964 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62096 2220 62160
rect 2284 62096 7740 62160
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62096 13740 62160
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62096 14220 62160
rect 14284 62096 19740 62160
rect 19804 62096 19820 62160
rect 19884 62096 19900 62160
rect 19964 62096 19980 62160
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62096 25740 62160
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62096 31740 62160
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62096 37740 62160
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62096 43740 62160
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62096 49740 62160
rect 49804 62096 49820 62160
rect 49884 62096 49900 62160
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62096 55740 62160
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62096 61740 62160
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62096 67740 62160
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62156 73740 62160
rect 68284 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 73740 62156
rect 68284 62096 73740 62100
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 75028 62160
rect 964 62080 75028 62096
rect 964 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62016 2220 62080
rect 2284 62016 7740 62080
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62016 13740 62080
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62016 14220 62080
rect 14284 62016 19740 62080
rect 19804 62016 19820 62080
rect 19884 62016 19900 62080
rect 19964 62016 19980 62080
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62016 25740 62080
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62016 31740 62080
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62016 37740 62080
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62016 43740 62080
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62016 49740 62080
rect 49804 62016 49820 62080
rect 49884 62016 49900 62080
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62016 55740 62080
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62016 61740 62080
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62016 67740 62080
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62076 73740 62080
rect 68284 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 73740 62076
rect 68284 62016 73740 62020
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 75028 62080
rect 964 62000 75028 62016
rect 964 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61936 2220 62000
rect 2284 61936 7740 62000
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61936 13740 62000
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61936 14220 62000
rect 14284 61936 19740 62000
rect 19804 61936 19820 62000
rect 19884 61936 19900 62000
rect 19964 61936 19980 62000
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61936 25740 62000
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61936 31740 62000
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61936 37740 62000
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61936 43740 62000
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61936 49740 62000
rect 49804 61936 49820 62000
rect 49884 61936 49900 62000
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61936 55740 62000
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61936 61740 62000
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61936 67740 62000
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61996 73740 62000
rect 68284 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 73740 61996
rect 68284 61936 73740 61940
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 75028 62000
rect 964 61912 75028 61936
rect 964 54592 75028 54616
rect 964 54528 4740 54592
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54528 10740 54592
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54528 16740 54592
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54528 17140 54592
rect 17204 54528 17220 54592
rect 17284 54528 22740 54592
rect 22804 54528 22820 54592
rect 22884 54528 22900 54592
rect 22964 54528 22980 54592
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54528 28740 54592
rect 28804 54528 28820 54592
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54528 34740 54592
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54528 40740 54592
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54528 46740 54592
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54528 52740 54592
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54528 58740 54592
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54528 59060 54592
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54588 64740 54592
rect 59284 54532 64216 54588
rect 64272 54532 64296 54588
rect 64352 54532 64376 54588
rect 64432 54532 64456 54588
rect 64512 54532 64740 54588
rect 59284 54528 64740 54532
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54588 75028 54592
rect 71284 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 75028 54588
rect 71284 54528 75028 54532
rect 964 54512 75028 54528
rect 964 54448 4740 54512
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54448 10740 54512
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54448 16740 54512
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54448 17140 54512
rect 17204 54448 17220 54512
rect 17284 54448 22740 54512
rect 22804 54448 22820 54512
rect 22884 54448 22900 54512
rect 22964 54448 22980 54512
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54448 28740 54512
rect 28804 54448 28820 54512
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54448 34740 54512
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54448 40740 54512
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54448 46740 54512
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54448 52740 54512
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54448 58740 54512
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54448 59060 54512
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54508 64740 54512
rect 59284 54452 64216 54508
rect 64272 54452 64296 54508
rect 64352 54452 64376 54508
rect 64432 54452 64456 54508
rect 64512 54452 64740 54508
rect 59284 54448 64740 54452
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54508 75028 54512
rect 71284 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 75028 54508
rect 71284 54448 75028 54452
rect 964 54432 75028 54448
rect 964 54368 4740 54432
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54368 10740 54432
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54368 16740 54432
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54368 17140 54432
rect 17204 54368 17220 54432
rect 17284 54368 22740 54432
rect 22804 54368 22820 54432
rect 22884 54368 22900 54432
rect 22964 54368 22980 54432
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54368 28740 54432
rect 28804 54368 28820 54432
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54368 34740 54432
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54368 40740 54432
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54368 46740 54432
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54368 52740 54432
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54368 58740 54432
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54368 59060 54432
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54428 64740 54432
rect 59284 54372 64216 54428
rect 64272 54372 64296 54428
rect 64352 54372 64376 54428
rect 64432 54372 64456 54428
rect 64512 54372 64740 54428
rect 59284 54368 64740 54372
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54428 75028 54432
rect 71284 54372 74216 54428
rect 74272 54372 74296 54428
rect 74352 54372 74376 54428
rect 74432 54372 74456 54428
rect 74512 54372 75028 54428
rect 71284 54368 75028 54372
rect 964 54352 75028 54368
rect 964 54288 4740 54352
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54288 10740 54352
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54288 16740 54352
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54288 17140 54352
rect 17204 54288 17220 54352
rect 17284 54288 22740 54352
rect 22804 54288 22820 54352
rect 22884 54288 22900 54352
rect 22964 54288 22980 54352
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54288 28740 54352
rect 28804 54288 28820 54352
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54288 34740 54352
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54288 40740 54352
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54288 46740 54352
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54288 52740 54352
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54288 58740 54352
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54288 59060 54352
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54348 64740 54352
rect 59284 54292 64216 54348
rect 64272 54292 64296 54348
rect 64352 54292 64376 54348
rect 64432 54292 64456 54348
rect 64512 54292 64740 54348
rect 59284 54288 64740 54292
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54348 75028 54352
rect 71284 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 75028 54348
rect 71284 54288 75028 54292
rect 964 54264 75028 54288
rect 63493 52594 63559 52597
rect 64086 52594 64092 52596
rect 63493 52592 64092 52594
rect 63493 52536 63498 52592
rect 63554 52536 64092 52592
rect 63493 52534 64092 52536
rect 63493 52531 63559 52534
rect 64086 52532 64092 52534
rect 64156 52532 64162 52596
rect 964 52240 75028 52264
rect 964 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52176 2220 52240
rect 2284 52176 7740 52240
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52176 13740 52240
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52176 14220 52240
rect 14284 52176 19740 52240
rect 19804 52176 19820 52240
rect 19884 52176 19900 52240
rect 19964 52176 19980 52240
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52176 25740 52240
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52176 31740 52240
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52176 37740 52240
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52176 43740 52240
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52176 49740 52240
rect 49804 52176 49820 52240
rect 49884 52176 49900 52240
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52176 55740 52240
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52176 61740 52240
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52176 67740 52240
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52236 73740 52240
rect 68284 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 73740 52236
rect 68284 52176 73740 52180
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 75028 52240
rect 964 52160 75028 52176
rect 964 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52096 2220 52160
rect 2284 52096 7740 52160
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52096 13740 52160
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52096 14220 52160
rect 14284 52096 19740 52160
rect 19804 52096 19820 52160
rect 19884 52096 19900 52160
rect 19964 52096 19980 52160
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52096 25740 52160
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52096 31740 52160
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52096 37740 52160
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52096 43740 52160
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52096 49740 52160
rect 49804 52096 49820 52160
rect 49884 52096 49900 52160
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52096 55740 52160
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52096 61740 52160
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52096 67740 52160
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52156 73740 52160
rect 68284 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 73740 52156
rect 68284 52096 73740 52100
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 75028 52160
rect 964 52080 75028 52096
rect 964 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52016 2220 52080
rect 2284 52016 7740 52080
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52016 13740 52080
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52016 14220 52080
rect 14284 52016 19740 52080
rect 19804 52016 19820 52080
rect 19884 52016 19900 52080
rect 19964 52016 19980 52080
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52016 25740 52080
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52016 31740 52080
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52016 37740 52080
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52016 43740 52080
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52016 49740 52080
rect 49804 52016 49820 52080
rect 49884 52016 49900 52080
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52016 55740 52080
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52016 61740 52080
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52016 67740 52080
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52076 73740 52080
rect 68284 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 73740 52076
rect 68284 52016 73740 52020
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 75028 52080
rect 964 52000 75028 52016
rect 964 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51936 2220 52000
rect 2284 51936 7740 52000
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51936 13740 52000
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51936 14220 52000
rect 14284 51936 19740 52000
rect 19804 51936 19820 52000
rect 19884 51936 19900 52000
rect 19964 51936 19980 52000
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51936 25740 52000
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51936 31740 52000
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51936 37740 52000
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51936 43740 52000
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51936 49740 52000
rect 49804 51936 49820 52000
rect 49884 51936 49900 52000
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51936 55740 52000
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51936 61740 52000
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51936 67740 52000
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51996 73740 52000
rect 68284 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 73740 51996
rect 68284 51936 73740 51940
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 75028 52000
rect 964 51912 75028 51936
rect 63493 50282 63559 50285
rect 64270 50282 64276 50284
rect 63493 50280 64276 50282
rect 63493 50224 63498 50280
rect 63554 50224 64276 50280
rect 63493 50222 64276 50224
rect 63493 50219 63559 50222
rect 64270 50220 64276 50222
rect 64340 50220 64346 50284
rect 62982 48724 62988 48788
rect 63052 48786 63058 48788
rect 63401 48786 63467 48789
rect 63052 48784 63467 48786
rect 63052 48728 63406 48784
rect 63462 48728 63467 48784
rect 63052 48726 63467 48728
rect 63052 48724 63058 48726
rect 63401 48723 63467 48726
rect 63493 48106 63559 48109
rect 64454 48106 64460 48108
rect 63493 48104 64460 48106
rect 63493 48048 63498 48104
rect 63554 48048 64460 48104
rect 63493 48046 64460 48048
rect 63493 48043 63559 48046
rect 64454 48044 64460 48046
rect 64524 48044 64530 48108
rect 63861 47700 63927 47701
rect 63861 47696 63908 47700
rect 63972 47698 63978 47700
rect 63861 47640 63866 47696
rect 63861 47636 63908 47640
rect 63972 47638 64018 47698
rect 63972 47636 63978 47638
rect 63861 47635 63927 47636
rect 964 44592 75028 44616
rect 964 44528 4740 44592
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44528 10740 44592
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44528 16740 44592
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44528 17140 44592
rect 17204 44528 17220 44592
rect 17284 44528 22740 44592
rect 22804 44528 22820 44592
rect 22884 44528 22900 44592
rect 22964 44528 22980 44592
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44528 28740 44592
rect 28804 44528 28820 44592
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44528 34740 44592
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44528 40740 44592
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44528 46740 44592
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44528 52740 44592
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44528 58740 44592
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44528 59060 44592
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44588 64740 44592
rect 59284 44532 64216 44588
rect 64272 44532 64296 44588
rect 64352 44532 64376 44588
rect 64432 44532 64456 44588
rect 64512 44532 64740 44588
rect 59284 44528 64740 44532
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44588 75028 44592
rect 71284 44532 74216 44588
rect 74272 44532 74296 44588
rect 74352 44532 74376 44588
rect 74432 44532 74456 44588
rect 74512 44532 75028 44588
rect 71284 44528 75028 44532
rect 964 44512 75028 44528
rect 964 44448 4740 44512
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44448 10740 44512
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44448 16740 44512
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44448 17140 44512
rect 17204 44448 17220 44512
rect 17284 44448 22740 44512
rect 22804 44448 22820 44512
rect 22884 44448 22900 44512
rect 22964 44448 22980 44512
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44448 28740 44512
rect 28804 44448 28820 44512
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44448 34740 44512
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44448 40740 44512
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44448 46740 44512
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44448 52740 44512
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44448 58740 44512
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44448 59060 44512
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44508 64740 44512
rect 59284 44452 64216 44508
rect 64272 44452 64296 44508
rect 64352 44452 64376 44508
rect 64432 44452 64456 44508
rect 64512 44452 64740 44508
rect 59284 44448 64740 44452
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44508 75028 44512
rect 71284 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 75028 44508
rect 71284 44448 75028 44452
rect 964 44432 75028 44448
rect 964 44368 4740 44432
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44368 10740 44432
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44368 16740 44432
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44368 17140 44432
rect 17204 44368 17220 44432
rect 17284 44368 22740 44432
rect 22804 44368 22820 44432
rect 22884 44368 22900 44432
rect 22964 44368 22980 44432
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44368 28740 44432
rect 28804 44368 28820 44432
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44368 34740 44432
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44368 40740 44432
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44368 46740 44432
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44368 52740 44432
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44368 58740 44432
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44368 59060 44432
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44428 64740 44432
rect 59284 44372 64216 44428
rect 64272 44372 64296 44428
rect 64352 44372 64376 44428
rect 64432 44372 64456 44428
rect 64512 44372 64740 44428
rect 59284 44368 64740 44372
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44428 75028 44432
rect 71284 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 75028 44428
rect 71284 44368 75028 44372
rect 964 44352 75028 44368
rect 964 44288 4740 44352
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44288 10740 44352
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44288 16740 44352
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44288 17140 44352
rect 17204 44288 17220 44352
rect 17284 44288 22740 44352
rect 22804 44288 22820 44352
rect 22884 44288 22900 44352
rect 22964 44288 22980 44352
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44288 28740 44352
rect 28804 44288 28820 44352
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44288 34740 44352
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44288 40740 44352
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44288 46740 44352
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44288 52740 44352
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44288 58740 44352
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44288 59060 44352
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44348 64740 44352
rect 59284 44292 64216 44348
rect 64272 44292 64296 44348
rect 64352 44292 64376 44348
rect 64432 44292 64456 44348
rect 64512 44292 64740 44348
rect 59284 44288 64740 44292
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44348 75028 44352
rect 71284 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 75028 44348
rect 71284 44288 75028 44292
rect 964 44264 75028 44288
rect 964 42240 75028 42264
rect 964 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42176 2220 42240
rect 2284 42176 7740 42240
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42176 13740 42240
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42176 14220 42240
rect 14284 42176 19740 42240
rect 19804 42176 19820 42240
rect 19884 42176 19900 42240
rect 19964 42176 19980 42240
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42176 25740 42240
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42176 31740 42240
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42176 37740 42240
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42176 43740 42240
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42176 49740 42240
rect 49804 42176 49820 42240
rect 49884 42176 49900 42240
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42176 55740 42240
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42176 61740 42240
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42176 67740 42240
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42236 73740 42240
rect 68284 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 73740 42236
rect 68284 42176 73740 42180
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 75028 42240
rect 964 42160 75028 42176
rect 964 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42096 2220 42160
rect 2284 42096 7740 42160
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42096 13740 42160
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42096 14220 42160
rect 14284 42096 19740 42160
rect 19804 42096 19820 42160
rect 19884 42096 19900 42160
rect 19964 42096 19980 42160
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42096 25740 42160
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42096 31740 42160
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42096 37740 42160
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42096 43740 42160
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42096 49740 42160
rect 49804 42096 49820 42160
rect 49884 42096 49900 42160
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42096 55740 42160
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42096 61740 42160
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42096 67740 42160
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42156 73740 42160
rect 68284 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 73740 42156
rect 68284 42096 73740 42100
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 75028 42160
rect 964 42080 75028 42096
rect 964 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42016 2220 42080
rect 2284 42016 7740 42080
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42016 13740 42080
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42016 14220 42080
rect 14284 42016 19740 42080
rect 19804 42016 19820 42080
rect 19884 42016 19900 42080
rect 19964 42016 19980 42080
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42016 25740 42080
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42016 31740 42080
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42016 37740 42080
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42016 43740 42080
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42016 49740 42080
rect 49804 42016 49820 42080
rect 49884 42016 49900 42080
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42016 55740 42080
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42016 61740 42080
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42016 67740 42080
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42076 73740 42080
rect 68284 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 73740 42076
rect 68284 42016 73740 42020
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 75028 42080
rect 964 42000 75028 42016
rect 964 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41936 2220 42000
rect 2284 41936 7740 42000
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41936 13740 42000
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41936 14220 42000
rect 14284 41936 19740 42000
rect 19804 41936 19820 42000
rect 19884 41936 19900 42000
rect 19964 41936 19980 42000
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41936 25740 42000
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41936 31740 42000
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41936 37740 42000
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41936 43740 42000
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41936 49740 42000
rect 49804 41936 49820 42000
rect 49884 41936 49900 42000
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41936 55740 42000
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41936 61740 42000
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41936 67740 42000
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41996 73740 42000
rect 68284 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 73740 41996
rect 68284 41936 73740 41940
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 75028 42000
rect 964 41912 75028 41936
rect 64965 40898 65031 40901
rect 65558 40898 65564 40900
rect 64965 40896 65564 40898
rect 64965 40840 64970 40896
rect 65026 40840 65564 40896
rect 64965 40838 65564 40840
rect 64965 40835 65031 40838
rect 65558 40836 65564 40838
rect 65628 40836 65634 40900
rect 64965 38858 65031 38861
rect 65742 38858 65748 38860
rect 64965 38856 65748 38858
rect 64965 38800 64970 38856
rect 65026 38800 65748 38856
rect 64965 38798 65748 38800
rect 64965 38795 65031 38798
rect 65742 38796 65748 38798
rect 65812 38796 65818 38860
rect 65517 34778 65583 34781
rect 65926 34778 65932 34780
rect 65517 34776 65932 34778
rect 65517 34720 65522 34776
rect 65578 34720 65932 34776
rect 65517 34718 65932 34720
rect 65517 34715 65583 34718
rect 65926 34716 65932 34718
rect 65996 34716 66002 34780
rect 964 34592 75028 34616
rect 964 34528 4740 34592
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34528 10740 34592
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34528 16740 34592
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34528 17140 34592
rect 17204 34528 17220 34592
rect 17284 34528 22740 34592
rect 22804 34528 22820 34592
rect 22884 34528 22900 34592
rect 22964 34528 22980 34592
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34528 28740 34592
rect 28804 34528 28820 34592
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34528 34740 34592
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34528 40740 34592
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34528 46740 34592
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34528 52740 34592
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34528 58740 34592
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34528 59060 34592
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34588 64740 34592
rect 59284 34532 64216 34588
rect 64272 34532 64296 34588
rect 64352 34532 64376 34588
rect 64432 34532 64456 34588
rect 64512 34532 64740 34588
rect 59284 34528 64740 34532
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34588 75028 34592
rect 71284 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 75028 34588
rect 71284 34528 75028 34532
rect 964 34512 75028 34528
rect 964 34448 4740 34512
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34448 10740 34512
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34448 16740 34512
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34448 17140 34512
rect 17204 34448 17220 34512
rect 17284 34448 22740 34512
rect 22804 34448 22820 34512
rect 22884 34448 22900 34512
rect 22964 34448 22980 34512
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34448 28740 34512
rect 28804 34448 28820 34512
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34448 34740 34512
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34448 40740 34512
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34448 46740 34512
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34448 52740 34512
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34448 58740 34512
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34448 59060 34512
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34508 64740 34512
rect 59284 34452 64216 34508
rect 64272 34452 64296 34508
rect 64352 34452 64376 34508
rect 64432 34452 64456 34508
rect 64512 34452 64740 34508
rect 59284 34448 64740 34452
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34508 75028 34512
rect 71284 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 75028 34508
rect 71284 34448 75028 34452
rect 964 34432 75028 34448
rect 964 34368 4740 34432
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34368 10740 34432
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34368 16740 34432
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34368 17140 34432
rect 17204 34368 17220 34432
rect 17284 34368 22740 34432
rect 22804 34368 22820 34432
rect 22884 34368 22900 34432
rect 22964 34368 22980 34432
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34368 28740 34432
rect 28804 34368 28820 34432
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34368 34740 34432
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34368 40740 34432
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34368 46740 34432
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34368 52740 34432
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34368 58740 34432
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34368 59060 34432
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34428 64740 34432
rect 59284 34372 64216 34428
rect 64272 34372 64296 34428
rect 64352 34372 64376 34428
rect 64432 34372 64456 34428
rect 64512 34372 64740 34428
rect 59284 34368 64740 34372
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34428 75028 34432
rect 71284 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 75028 34428
rect 71284 34368 75028 34372
rect 964 34352 75028 34368
rect 964 34288 4740 34352
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34288 10740 34352
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34288 16740 34352
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34288 17140 34352
rect 17204 34288 17220 34352
rect 17284 34288 22740 34352
rect 22804 34288 22820 34352
rect 22884 34288 22900 34352
rect 22964 34288 22980 34352
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34288 28740 34352
rect 28804 34288 28820 34352
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34288 34740 34352
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34288 40740 34352
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34288 46740 34352
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34288 52740 34352
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34288 58740 34352
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34288 59060 34352
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34348 64740 34352
rect 59284 34292 64216 34348
rect 64272 34292 64296 34348
rect 64352 34292 64376 34348
rect 64432 34292 64456 34348
rect 64512 34292 64740 34348
rect 59284 34288 64740 34292
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34348 75028 34352
rect 71284 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 75028 34348
rect 71284 34288 75028 34292
rect 964 34264 75028 34288
rect 65609 33282 65675 33285
rect 68502 33282 68508 33284
rect 65609 33280 68508 33282
rect 65609 33224 65614 33280
rect 65670 33224 68508 33280
rect 65609 33222 68508 33224
rect 65609 33219 65675 33222
rect 68502 33220 68508 33222
rect 68572 33220 68578 33284
rect 964 32240 75028 32264
rect 964 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32176 2220 32240
rect 2284 32176 7740 32240
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32176 13740 32240
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32176 14220 32240
rect 14284 32176 19740 32240
rect 19804 32176 19820 32240
rect 19884 32176 19900 32240
rect 19964 32176 19980 32240
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32176 25740 32240
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32176 31740 32240
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32176 37740 32240
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32176 43740 32240
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32176 49740 32240
rect 49804 32176 49820 32240
rect 49884 32176 49900 32240
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32176 55740 32240
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32176 61740 32240
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32176 67740 32240
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32236 73740 32240
rect 68284 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 73740 32236
rect 68284 32176 73740 32180
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 75028 32240
rect 964 32160 75028 32176
rect 964 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32096 2220 32160
rect 2284 32096 7740 32160
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32096 13740 32160
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32096 14220 32160
rect 14284 32096 19740 32160
rect 19804 32096 19820 32160
rect 19884 32096 19900 32160
rect 19964 32096 19980 32160
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32096 25740 32160
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32096 31740 32160
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32096 37740 32160
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32096 43740 32160
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32096 49740 32160
rect 49804 32096 49820 32160
rect 49884 32096 49900 32160
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32096 55740 32160
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32096 61740 32160
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32096 67740 32160
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32156 73740 32160
rect 68284 32100 71864 32156
rect 71920 32100 71944 32156
rect 72000 32100 72024 32156
rect 72080 32100 72104 32156
rect 72160 32100 73740 32156
rect 68284 32096 73740 32100
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 75028 32160
rect 964 32080 75028 32096
rect 964 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32016 2220 32080
rect 2284 32016 7740 32080
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32016 13740 32080
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32016 14220 32080
rect 14284 32016 19740 32080
rect 19804 32016 19820 32080
rect 19884 32016 19900 32080
rect 19964 32016 19980 32080
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32016 25740 32080
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32016 31740 32080
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32016 37740 32080
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32016 43740 32080
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32016 49740 32080
rect 49804 32016 49820 32080
rect 49884 32016 49900 32080
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32016 55740 32080
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32016 61740 32080
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32016 67740 32080
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32076 73740 32080
rect 68284 32020 71864 32076
rect 71920 32020 71944 32076
rect 72000 32020 72024 32076
rect 72080 32020 72104 32076
rect 72160 32020 73740 32076
rect 68284 32016 73740 32020
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 75028 32080
rect 964 32000 75028 32016
rect 964 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31936 2220 32000
rect 2284 31936 7740 32000
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31936 13740 32000
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31936 14220 32000
rect 14284 31936 19740 32000
rect 19804 31936 19820 32000
rect 19884 31936 19900 32000
rect 19964 31936 19980 32000
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31936 25740 32000
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31936 31740 32000
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31936 37740 32000
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31936 43740 32000
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31936 49740 32000
rect 49804 31936 49820 32000
rect 49884 31936 49900 32000
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31936 55740 32000
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31936 61740 32000
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31936 67740 32000
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31996 73740 32000
rect 68284 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 73740 31996
rect 68284 31936 73740 31940
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 75028 32000
rect 964 31912 75028 31936
rect 67357 26484 67423 26485
rect 67357 26480 67404 26484
rect 67468 26482 67474 26484
rect 67357 26424 67362 26480
rect 67357 26420 67404 26424
rect 67468 26422 67514 26482
rect 67468 26420 67474 26422
rect 67357 26419 67423 26420
rect 63166 26148 63172 26212
rect 63236 26210 63242 26212
rect 63677 26210 63743 26213
rect 63236 26208 63743 26210
rect 63236 26152 63682 26208
rect 63738 26152 63743 26208
rect 63236 26150 63743 26152
rect 63236 26148 63242 26150
rect 63677 26147 63743 26150
rect 67398 26012 67404 26076
rect 67468 26074 67474 26076
rect 67541 26074 67607 26077
rect 67468 26072 67607 26074
rect 67468 26016 67546 26072
rect 67602 26016 67607 26072
rect 67468 26014 67607 26016
rect 67468 26012 67474 26014
rect 67541 26011 67607 26014
rect 964 24592 75028 24616
rect 964 24528 4740 24592
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24528 10740 24592
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24528 16740 24592
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24528 17140 24592
rect 17204 24528 17220 24592
rect 17284 24528 22740 24592
rect 22804 24528 22820 24592
rect 22884 24528 22900 24592
rect 22964 24528 22980 24592
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24528 28740 24592
rect 28804 24528 28820 24592
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24528 34740 24592
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24528 40740 24592
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24528 46740 24592
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24528 52740 24592
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24528 58740 24592
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24528 59060 24592
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24588 64740 24592
rect 59284 24532 64216 24588
rect 64272 24532 64296 24588
rect 64352 24532 64376 24588
rect 64432 24532 64456 24588
rect 64512 24532 64740 24588
rect 59284 24528 64740 24532
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24588 75028 24592
rect 71284 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 75028 24588
rect 71284 24528 75028 24532
rect 964 24512 75028 24528
rect 964 24448 4740 24512
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24448 10740 24512
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24448 16740 24512
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24448 17140 24512
rect 17204 24448 17220 24512
rect 17284 24448 22740 24512
rect 22804 24448 22820 24512
rect 22884 24448 22900 24512
rect 22964 24448 22980 24512
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24448 28740 24512
rect 28804 24448 28820 24512
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24448 34740 24512
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24448 40740 24512
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24448 46740 24512
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24448 52740 24512
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24448 58740 24512
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24448 59060 24512
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24508 64740 24512
rect 59284 24452 64216 24508
rect 64272 24452 64296 24508
rect 64352 24452 64376 24508
rect 64432 24452 64456 24508
rect 64512 24452 64740 24508
rect 59284 24448 64740 24452
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24508 75028 24512
rect 71284 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 75028 24508
rect 71284 24448 75028 24452
rect 964 24432 75028 24448
rect 964 24368 4740 24432
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24368 10740 24432
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24368 16740 24432
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24368 17140 24432
rect 17204 24368 17220 24432
rect 17284 24368 22740 24432
rect 22804 24368 22820 24432
rect 22884 24368 22900 24432
rect 22964 24368 22980 24432
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24368 28740 24432
rect 28804 24368 28820 24432
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24368 34740 24432
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24368 40740 24432
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24368 46740 24432
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24368 52740 24432
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24368 58740 24432
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24368 59060 24432
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24428 64740 24432
rect 59284 24372 64216 24428
rect 64272 24372 64296 24428
rect 64352 24372 64376 24428
rect 64432 24372 64456 24428
rect 64512 24372 64740 24428
rect 59284 24368 64740 24372
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24428 75028 24432
rect 71284 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 75028 24428
rect 71284 24368 75028 24372
rect 964 24352 75028 24368
rect 964 24288 4740 24352
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24288 10740 24352
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24288 16740 24352
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24288 17140 24352
rect 17204 24288 17220 24352
rect 17284 24288 22740 24352
rect 22804 24288 22820 24352
rect 22884 24288 22900 24352
rect 22964 24288 22980 24352
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24288 28740 24352
rect 28804 24288 28820 24352
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24288 34740 24352
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24288 40740 24352
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24288 46740 24352
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24288 52740 24352
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24288 58740 24352
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24288 59060 24352
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24348 64740 24352
rect 59284 24292 64216 24348
rect 64272 24292 64296 24348
rect 64352 24292 64376 24348
rect 64432 24292 64456 24348
rect 64512 24292 64740 24348
rect 59284 24288 64740 24292
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24348 75028 24352
rect 71284 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 75028 24348
rect 71284 24288 75028 24292
rect 964 24264 75028 24288
rect 66478 23564 66484 23628
rect 66548 23626 66554 23628
rect 67633 23626 67699 23629
rect 66548 23624 67699 23626
rect 66548 23568 67638 23624
rect 67694 23568 67699 23624
rect 66548 23566 67699 23568
rect 66548 23564 66554 23566
rect 67633 23563 67699 23566
rect 66294 23428 66300 23492
rect 66364 23490 66370 23492
rect 66437 23490 66503 23493
rect 66364 23488 66503 23490
rect 66364 23432 66442 23488
rect 66498 23432 66503 23488
rect 66364 23430 66503 23432
rect 66364 23428 66370 23430
rect 66437 23427 66503 23430
rect 66437 22402 66503 22405
rect 66662 22402 66668 22404
rect 66437 22400 66668 22402
rect 66437 22344 66442 22400
rect 66498 22344 66668 22400
rect 66437 22342 66668 22344
rect 66437 22339 66503 22342
rect 66662 22340 66668 22342
rect 66732 22340 66738 22404
rect 964 22240 75028 22264
rect 964 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22176 2220 22240
rect 2284 22176 7740 22240
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22176 13740 22240
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22176 14220 22240
rect 14284 22176 19740 22240
rect 19804 22176 19820 22240
rect 19884 22176 19900 22240
rect 19964 22176 19980 22240
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22176 25740 22240
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22176 31740 22240
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22176 37740 22240
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22176 43740 22240
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22176 49740 22240
rect 49804 22176 49820 22240
rect 49884 22176 49900 22240
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22176 55740 22240
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22176 61740 22240
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22176 67740 22240
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22236 73740 22240
rect 68284 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 73740 22236
rect 68284 22176 73740 22180
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 75028 22240
rect 964 22160 75028 22176
rect 964 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22096 2220 22160
rect 2284 22096 7740 22160
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22096 13740 22160
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22096 14220 22160
rect 14284 22096 19740 22160
rect 19804 22096 19820 22160
rect 19884 22096 19900 22160
rect 19964 22096 19980 22160
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22096 25740 22160
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22096 31740 22160
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22096 37740 22160
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22096 43740 22160
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22096 49740 22160
rect 49804 22096 49820 22160
rect 49884 22096 49900 22160
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22096 55740 22160
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22096 61740 22160
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22096 67740 22160
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22156 73740 22160
rect 68284 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 73740 22156
rect 68284 22096 73740 22100
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 75028 22160
rect 964 22080 75028 22096
rect 964 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22016 2220 22080
rect 2284 22016 7740 22080
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22016 13740 22080
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22016 14220 22080
rect 14284 22016 19740 22080
rect 19804 22016 19820 22080
rect 19884 22016 19900 22080
rect 19964 22016 19980 22080
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22016 25740 22080
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22016 31740 22080
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22016 37740 22080
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22016 43740 22080
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22016 49740 22080
rect 49804 22016 49820 22080
rect 49884 22016 49900 22080
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22016 55740 22080
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22016 61740 22080
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22016 67740 22080
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22076 73740 22080
rect 68284 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 73740 22076
rect 68284 22016 73740 22020
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 75028 22080
rect 964 22000 75028 22016
rect 964 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21936 2220 22000
rect 2284 21936 7740 22000
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21936 13740 22000
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21936 14220 22000
rect 14284 21936 19740 22000
rect 19804 21936 19820 22000
rect 19884 21936 19900 22000
rect 19964 21936 19980 22000
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21936 25740 22000
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21936 31740 22000
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21936 37740 22000
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21936 43740 22000
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21936 49740 22000
rect 49804 21936 49820 22000
rect 49884 21936 49900 22000
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21936 55740 22000
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21936 61740 22000
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21936 67740 22000
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21996 73740 22000
rect 68284 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 73740 21996
rect 68284 21936 73740 21940
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 75028 22000
rect 964 21912 75028 21936
rect 63534 16492 63540 16556
rect 63604 16554 63610 16556
rect 63769 16554 63835 16557
rect 63604 16552 63835 16554
rect 63604 16496 63774 16552
rect 63830 16496 63835 16552
rect 63604 16494 63835 16496
rect 63604 16492 63610 16494
rect 63769 16491 63835 16494
rect 63718 14724 63724 14788
rect 63788 14786 63794 14788
rect 64454 14786 64460 14788
rect 63788 14726 64460 14786
rect 63788 14724 63794 14726
rect 64454 14724 64460 14726
rect 64524 14724 64530 14788
rect 964 14592 75028 14616
rect 964 14528 4740 14592
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14528 10740 14592
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14528 16740 14592
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14528 17140 14592
rect 17204 14528 17220 14592
rect 17284 14528 22740 14592
rect 22804 14528 22820 14592
rect 22884 14528 22900 14592
rect 22964 14528 22980 14592
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14528 28740 14592
rect 28804 14528 28820 14592
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14528 34740 14592
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14528 40740 14592
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14528 46740 14592
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14528 52740 14592
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14528 58740 14592
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14528 59060 14592
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14588 64740 14592
rect 59284 14532 64216 14588
rect 64272 14532 64296 14588
rect 64352 14532 64376 14588
rect 64432 14532 64456 14588
rect 64512 14532 64740 14588
rect 59284 14528 64740 14532
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14588 75028 14592
rect 71284 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 75028 14588
rect 71284 14528 75028 14532
rect 964 14512 75028 14528
rect 964 14448 4740 14512
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14448 10740 14512
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14448 16740 14512
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14448 17140 14512
rect 17204 14448 17220 14512
rect 17284 14448 22740 14512
rect 22804 14448 22820 14512
rect 22884 14448 22900 14512
rect 22964 14448 22980 14512
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14448 28740 14512
rect 28804 14448 28820 14512
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14448 34740 14512
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14448 40740 14512
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14448 46740 14512
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14448 52740 14512
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14448 58740 14512
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14448 59060 14512
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14508 64740 14512
rect 59284 14452 64216 14508
rect 64272 14452 64296 14508
rect 64352 14452 64376 14508
rect 64432 14452 64456 14508
rect 64512 14452 64740 14508
rect 59284 14448 64740 14452
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14508 75028 14512
rect 71284 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 75028 14508
rect 71284 14448 75028 14452
rect 964 14432 75028 14448
rect 964 14368 4740 14432
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14368 10740 14432
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14368 16740 14432
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14368 17140 14432
rect 17204 14368 17220 14432
rect 17284 14368 22740 14432
rect 22804 14368 22820 14432
rect 22884 14368 22900 14432
rect 22964 14368 22980 14432
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14368 28740 14432
rect 28804 14368 28820 14432
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14368 34740 14432
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14368 40740 14432
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14368 46740 14432
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14368 52740 14432
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14368 58740 14432
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14368 59060 14432
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14428 64740 14432
rect 59284 14372 64216 14428
rect 64272 14372 64296 14428
rect 64352 14372 64376 14428
rect 64432 14372 64456 14428
rect 64512 14372 64740 14428
rect 59284 14368 64740 14372
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14428 75028 14432
rect 71284 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 75028 14428
rect 71284 14368 75028 14372
rect 964 14352 75028 14368
rect 964 14288 4740 14352
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14288 10740 14352
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14288 16740 14352
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14288 17140 14352
rect 17204 14288 17220 14352
rect 17284 14288 22740 14352
rect 22804 14288 22820 14352
rect 22884 14288 22900 14352
rect 22964 14288 22980 14352
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14288 28740 14352
rect 28804 14288 28820 14352
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14288 34740 14352
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14288 40740 14352
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14288 46740 14352
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14288 52740 14352
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14288 58740 14352
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14288 59060 14352
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14348 64740 14352
rect 59284 14292 64216 14348
rect 64272 14292 64296 14348
rect 64352 14292 64376 14348
rect 64432 14292 64456 14348
rect 64512 14292 64740 14348
rect 59284 14288 64740 14292
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14348 75028 14352
rect 71284 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 75028 14348
rect 71284 14288 75028 14292
rect 964 14264 75028 14288
rect 64873 12746 64939 12749
rect 66846 12746 66852 12748
rect 64873 12744 66852 12746
rect 64873 12688 64878 12744
rect 64934 12688 66852 12744
rect 64873 12686 66852 12688
rect 64873 12683 64939 12686
rect 66846 12684 66852 12686
rect 66916 12684 66922 12748
rect 64086 12548 64092 12612
rect 64156 12610 64162 12612
rect 64873 12610 64939 12613
rect 64156 12608 64939 12610
rect 64156 12552 64878 12608
rect 64934 12552 64939 12608
rect 64156 12550 64939 12552
rect 64156 12548 64162 12550
rect 64873 12547 64939 12550
rect 964 12240 75028 12264
rect 964 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12176 2220 12240
rect 2284 12176 7740 12240
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12176 13740 12240
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12176 14220 12240
rect 14284 12176 19740 12240
rect 19804 12176 19820 12240
rect 19884 12176 19900 12240
rect 19964 12176 19980 12240
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12176 25740 12240
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12176 31740 12240
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12176 37740 12240
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12176 43740 12240
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12176 49740 12240
rect 49804 12176 49820 12240
rect 49884 12176 49900 12240
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12176 55740 12240
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12176 61740 12240
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12176 67740 12240
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12236 73740 12240
rect 68284 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 73740 12236
rect 68284 12176 73740 12180
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 75028 12240
rect 964 12160 75028 12176
rect 964 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12096 2220 12160
rect 2284 12096 7740 12160
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12096 13740 12160
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12096 14220 12160
rect 14284 12096 19740 12160
rect 19804 12096 19820 12160
rect 19884 12096 19900 12160
rect 19964 12096 19980 12160
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12096 25740 12160
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12096 31740 12160
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12096 37740 12160
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12096 43740 12160
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12096 49740 12160
rect 49804 12096 49820 12160
rect 49884 12096 49900 12160
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12096 55740 12160
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12096 61740 12160
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12096 67740 12160
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12156 73740 12160
rect 68284 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 73740 12156
rect 68284 12096 73740 12100
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 75028 12160
rect 964 12080 75028 12096
rect 964 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12016 2220 12080
rect 2284 12016 7740 12080
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12016 13740 12080
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12016 14220 12080
rect 14284 12016 19740 12080
rect 19804 12016 19820 12080
rect 19884 12016 19900 12080
rect 19964 12016 19980 12080
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12016 25740 12080
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12016 31740 12080
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12016 37740 12080
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12016 43740 12080
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12016 49740 12080
rect 49804 12016 49820 12080
rect 49884 12016 49900 12080
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12016 55740 12080
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12016 61740 12080
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12016 67740 12080
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12076 73740 12080
rect 68284 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 73740 12076
rect 68284 12016 73740 12020
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 75028 12080
rect 964 12000 75028 12016
rect 964 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2220 12000
rect 2284 11936 7740 12000
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11936 13740 12000
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11936 14220 12000
rect 14284 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11936 25740 12000
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11936 31740 12000
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 37740 12000
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11936 43740 12000
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11936 49740 12000
rect 49804 11936 49820 12000
rect 49884 11936 49900 12000
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11936 55740 12000
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11936 61740 12000
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11936 67740 12000
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11996 73740 12000
rect 68284 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 73740 11996
rect 68284 11936 73740 11940
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 75028 12000
rect 964 11912 75028 11936
rect 63493 11796 63559 11797
rect 63493 11794 63540 11796
rect 63448 11792 63540 11794
rect 63448 11736 63498 11792
rect 63448 11734 63540 11736
rect 63493 11732 63540 11734
rect 63604 11732 63610 11796
rect 64270 11732 64276 11796
rect 64340 11794 64346 11796
rect 64873 11794 64939 11797
rect 64340 11792 64939 11794
rect 64340 11736 64878 11792
rect 64934 11736 64939 11792
rect 64340 11734 64939 11736
rect 64340 11732 64346 11734
rect 63493 11731 63559 11732
rect 64873 11731 64939 11734
rect 63350 11596 63356 11660
rect 63420 11658 63426 11660
rect 63902 11658 63908 11660
rect 63420 11598 63908 11658
rect 63420 11596 63426 11598
rect 63902 11596 63908 11598
rect 63972 11596 63978 11660
rect 64045 11250 64111 11253
rect 64045 11248 64154 11250
rect 64045 11192 64050 11248
rect 64106 11192 64154 11248
rect 64045 11187 64154 11192
rect 64094 11116 64154 11187
rect 64086 11052 64092 11116
rect 64156 11052 64162 11116
rect 63401 10708 63467 10709
rect 63350 10706 63356 10708
rect 63310 10646 63356 10706
rect 63420 10704 63467 10708
rect 63462 10648 63467 10704
rect 63350 10644 63356 10646
rect 63420 10644 63467 10648
rect 63401 10643 63467 10644
rect 64045 7986 64111 7989
rect 63726 7984 64111 7986
rect 63726 7928 64050 7984
rect 64106 7928 64111 7984
rect 63726 7926 64111 7928
rect 59553 7850 59619 7853
rect 63726 7850 63786 7926
rect 64045 7923 64111 7926
rect 59553 7848 63786 7850
rect 59553 7792 59558 7848
rect 59614 7792 63786 7848
rect 59553 7790 63786 7792
rect 59553 7787 59619 7790
rect 41045 7714 41111 7717
rect 63902 7714 63908 7716
rect 41045 7712 63908 7714
rect 41045 7656 41050 7712
rect 41106 7656 63908 7712
rect 41045 7654 63908 7656
rect 41045 7651 41111 7654
rect 63902 7652 63908 7654
rect 63972 7652 63978 7716
rect 34053 7578 34119 7581
rect 62982 7578 62988 7580
rect 34053 7576 62988 7578
rect 34053 7520 34058 7576
rect 34114 7520 62988 7576
rect 34053 7518 62988 7520
rect 34053 7515 34119 7518
rect 62982 7516 62988 7518
rect 63052 7516 63058 7580
rect 59169 7442 59235 7445
rect 67173 7442 67239 7445
rect 59169 7440 67239 7442
rect 59169 7384 59174 7440
rect 59230 7384 67178 7440
rect 67234 7384 67239 7440
rect 59169 7382 67239 7384
rect 59169 7379 59235 7382
rect 67173 7379 67239 7382
rect 63350 7244 63356 7308
rect 63420 7306 63426 7308
rect 63493 7306 63559 7309
rect 63420 7304 63559 7306
rect 63420 7248 63498 7304
rect 63554 7248 63559 7304
rect 63420 7246 63559 7248
rect 63420 7244 63426 7246
rect 63493 7243 63559 7246
rect 59629 7034 59695 7037
rect 64086 7034 64092 7036
rect 59629 7032 64092 7034
rect 59629 6976 59634 7032
rect 59690 6976 64092 7032
rect 59629 6974 64092 6976
rect 59629 6971 59695 6974
rect 64086 6972 64092 6974
rect 64156 6972 64162 7036
rect 30281 6898 30347 6901
rect 30281 6896 60750 6898
rect 30281 6840 30286 6896
rect 30342 6840 60750 6896
rect 30281 6838 60750 6840
rect 30281 6835 30347 6838
rect 29637 6762 29703 6765
rect 60690 6762 60750 6838
rect 65558 6762 65564 6764
rect 29637 6760 51090 6762
rect 29637 6704 29642 6760
rect 29698 6704 51090 6760
rect 29637 6702 51090 6704
rect 60690 6702 65564 6762
rect 29637 6699 29703 6702
rect 29269 6626 29335 6629
rect 51030 6626 51090 6702
rect 65558 6700 65564 6702
rect 65628 6700 65634 6764
rect 65742 6626 65748 6628
rect 29269 6624 41430 6626
rect 29269 6568 29274 6624
rect 29330 6568 41430 6624
rect 29269 6566 41430 6568
rect 51030 6566 65748 6626
rect 29269 6563 29335 6566
rect 41370 6490 41430 6566
rect 65742 6564 65748 6566
rect 65812 6564 65818 6628
rect 66069 6490 66135 6493
rect 41370 6488 66135 6490
rect 41370 6432 66074 6488
rect 66130 6432 66135 6488
rect 41370 6430 66135 6432
rect 66069 6427 66135 6430
rect 56501 6354 56567 6357
rect 63585 6354 63651 6357
rect 56501 6352 63651 6354
rect 56501 6296 56506 6352
rect 56562 6296 63590 6352
rect 63646 6296 63651 6352
rect 56501 6294 63651 6296
rect 56501 6291 56567 6294
rect 63585 6291 63651 6294
rect 64873 6354 64939 6357
rect 66478 6354 66484 6356
rect 64873 6352 66484 6354
rect 64873 6296 64878 6352
rect 64934 6296 66484 6352
rect 64873 6294 66484 6296
rect 64873 6291 64939 6294
rect 66478 6292 66484 6294
rect 66548 6292 66554 6356
rect 55765 6218 55831 6221
rect 66846 6218 66852 6220
rect 55765 6216 66852 6218
rect 55765 6160 55770 6216
rect 55826 6160 66852 6216
rect 55765 6158 66852 6160
rect 55765 6155 55831 6158
rect 66846 6156 66852 6158
rect 66916 6156 66922 6220
rect 49509 6082 49575 6085
rect 57513 6082 57579 6085
rect 49509 6080 57579 6082
rect 49509 6024 49514 6080
rect 49570 6024 57518 6080
rect 57574 6024 57579 6080
rect 49509 6022 57579 6024
rect 49509 6019 49575 6022
rect 57513 6019 57579 6022
rect 58157 6082 58223 6085
rect 62757 6082 62823 6085
rect 58157 6080 62823 6082
rect 58157 6024 58162 6080
rect 58218 6024 62762 6080
rect 62818 6024 62823 6080
rect 58157 6022 62823 6024
rect 58157 6019 58223 6022
rect 62757 6019 62823 6022
rect 63125 6082 63191 6085
rect 65926 6082 65932 6084
rect 63125 6080 65932 6082
rect 63125 6024 63130 6080
rect 63186 6024 65932 6080
rect 63125 6022 65932 6024
rect 63125 6019 63191 6022
rect 65926 6020 65932 6022
rect 65996 6020 66002 6084
rect 25865 5946 25931 5949
rect 44633 5946 44699 5949
rect 64781 5946 64847 5949
rect 25865 5944 41430 5946
rect 25865 5888 25870 5944
rect 25926 5888 41430 5944
rect 25865 5886 41430 5888
rect 25865 5883 25931 5886
rect 39982 5748 39988 5812
rect 40052 5810 40058 5812
rect 40401 5810 40467 5813
rect 40052 5808 40467 5810
rect 40052 5752 40406 5808
rect 40462 5752 40467 5808
rect 40052 5750 40467 5752
rect 41370 5810 41430 5886
rect 44633 5944 64847 5946
rect 44633 5888 44638 5944
rect 44694 5888 64786 5944
rect 64842 5888 64847 5944
rect 44633 5886 64847 5888
rect 44633 5883 44699 5886
rect 64781 5883 64847 5886
rect 55765 5810 55831 5813
rect 41370 5808 55831 5810
rect 41370 5752 55770 5808
rect 55826 5752 55831 5808
rect 41370 5750 55831 5752
rect 40052 5748 40058 5750
rect 40401 5747 40467 5750
rect 55765 5747 55831 5750
rect 62941 5810 63007 5813
rect 63166 5810 63172 5812
rect 62941 5808 63172 5810
rect 62941 5752 62946 5808
rect 63002 5752 63172 5808
rect 62941 5750 63172 5752
rect 62941 5747 63007 5750
rect 63166 5748 63172 5750
rect 63236 5748 63242 5812
rect 63401 5810 63467 5813
rect 69013 5810 69079 5813
rect 63401 5808 69079 5810
rect 63401 5752 63406 5808
rect 63462 5752 69018 5808
rect 69074 5752 69079 5808
rect 63401 5750 69079 5752
rect 63401 5747 63467 5750
rect 69013 5747 69079 5750
rect 36997 5674 37063 5677
rect 41689 5674 41755 5677
rect 68502 5674 68508 5676
rect 36997 5672 68508 5674
rect 36997 5616 37002 5672
rect 37058 5616 41694 5672
rect 41750 5616 68508 5672
rect 36997 5614 68508 5616
rect 36997 5611 37063 5614
rect 41689 5611 41755 5614
rect 68502 5612 68508 5614
rect 68572 5612 68578 5676
rect 46013 5538 46079 5541
rect 55857 5538 55923 5541
rect 46013 5536 55923 5538
rect 46013 5480 46018 5536
rect 46074 5480 55862 5536
rect 55918 5480 55923 5536
rect 46013 5478 55923 5480
rect 46013 5475 46079 5478
rect 55857 5475 55923 5478
rect 60917 5538 60983 5541
rect 64965 5538 65031 5541
rect 60917 5536 65031 5538
rect 60917 5480 60922 5536
rect 60978 5480 64970 5536
rect 65026 5480 65031 5536
rect 60917 5478 65031 5480
rect 60917 5475 60983 5478
rect 64965 5475 65031 5478
rect 28441 5402 28507 5405
rect 63125 5402 63191 5405
rect 28441 5400 63191 5402
rect 28441 5344 28446 5400
rect 28502 5344 63130 5400
rect 63186 5344 63191 5400
rect 28441 5342 63191 5344
rect 28441 5339 28507 5342
rect 63125 5339 63191 5342
rect 63401 5402 63467 5405
rect 69105 5402 69171 5405
rect 63401 5400 69171 5402
rect 63401 5344 63406 5400
rect 63462 5344 69110 5400
rect 69166 5344 69171 5400
rect 63401 5342 69171 5344
rect 63401 5339 63467 5342
rect 69105 5339 69171 5342
rect 30833 5266 30899 5269
rect 70485 5266 70551 5269
rect 30833 5264 70551 5266
rect 30833 5208 30838 5264
rect 30894 5208 70490 5264
rect 70546 5208 70551 5264
rect 30833 5206 70551 5208
rect 30833 5203 30899 5206
rect 70485 5203 70551 5206
rect 25865 5130 25931 5133
rect 30373 5130 30439 5133
rect 25865 5128 30439 5130
rect 25865 5072 25870 5128
rect 25926 5072 30378 5128
rect 30434 5072 30439 5128
rect 25865 5070 30439 5072
rect 25865 5067 25931 5070
rect 30373 5067 30439 5070
rect 44081 5130 44147 5133
rect 47577 5130 47643 5133
rect 44081 5128 47643 5130
rect 44081 5072 44086 5128
rect 44142 5072 47582 5128
rect 47638 5072 47643 5128
rect 44081 5070 47643 5072
rect 44081 5067 44147 5070
rect 47577 5067 47643 5070
rect 55857 5130 55923 5133
rect 64270 5130 64276 5132
rect 55857 5128 64276 5130
rect 55857 5072 55862 5128
rect 55918 5072 64276 5128
rect 55857 5070 64276 5072
rect 55857 5067 55923 5070
rect 64270 5068 64276 5070
rect 64340 5068 64346 5132
rect 28993 4994 29059 4997
rect 29637 4994 29703 4997
rect 28993 4992 29703 4994
rect 28993 4936 28998 4992
rect 29054 4936 29642 4992
rect 29698 4936 29703 4992
rect 28993 4934 29703 4936
rect 28993 4931 29059 4934
rect 29637 4931 29703 4934
rect 44725 4994 44791 4997
rect 64454 4994 64460 4996
rect 44725 4992 64460 4994
rect 44725 4936 44730 4992
rect 44786 4936 64460 4992
rect 44725 4934 64460 4936
rect 44725 4931 44791 4934
rect 64454 4932 64460 4934
rect 64524 4932 64530 4996
rect 46657 4858 46723 4861
rect 63401 4858 63467 4861
rect 46657 4856 63467 4858
rect 46657 4800 46662 4856
rect 46718 4800 63406 4856
rect 63462 4800 63467 4856
rect 46657 4798 63467 4800
rect 46657 4795 46723 4798
rect 63401 4795 63467 4798
rect 63585 4858 63651 4861
rect 66662 4858 66668 4860
rect 63585 4856 66668 4858
rect 63585 4800 63590 4856
rect 63646 4800 66668 4856
rect 63585 4798 66668 4800
rect 63585 4795 63651 4798
rect 66662 4796 66668 4798
rect 66732 4796 66738 4860
rect 964 4592 75028 4616
rect 964 4588 4740 4592
rect 964 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4740 4588
rect 964 4528 4740 4532
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4588 16740 4592
rect 11284 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 16740 4588
rect 11284 4528 16740 4532
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4588 28740 4592
rect 23284 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 28740 4588
rect 23284 4528 28740 4532
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4588 34740 4592
rect 29284 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34740 4588
rect 29284 4528 34740 4532
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4588 46740 4592
rect 41284 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 46740 4588
rect 41284 4528 46740 4532
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4588 58740 4592
rect 53284 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 58740 4588
rect 53284 4528 58740 4532
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4588 64740 4592
rect 59284 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64740 4588
rect 59284 4528 64740 4532
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4588 75028 4592
rect 71284 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 75028 4588
rect 71284 4528 75028 4532
rect 964 4512 75028 4528
rect 964 4508 4740 4512
rect 964 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4740 4508
rect 964 4448 4740 4452
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4508 16740 4512
rect 11284 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 16740 4508
rect 11284 4448 16740 4452
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4508 28740 4512
rect 23284 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 28740 4508
rect 23284 4448 28740 4452
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4508 34740 4512
rect 29284 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34740 4508
rect 29284 4448 34740 4452
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4508 46740 4512
rect 41284 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 46740 4508
rect 41284 4448 46740 4452
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4508 58740 4512
rect 53284 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 58740 4508
rect 53284 4448 58740 4452
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4508 64740 4512
rect 59284 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64740 4508
rect 59284 4448 64740 4452
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4508 75028 4512
rect 71284 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 75028 4508
rect 71284 4448 75028 4452
rect 964 4432 75028 4448
rect 964 4428 4740 4432
rect 964 4372 4216 4428
rect 4272 4372 4296 4428
rect 4352 4372 4376 4428
rect 4432 4372 4456 4428
rect 4512 4372 4740 4428
rect 964 4368 4740 4372
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4428 16740 4432
rect 11284 4372 14216 4428
rect 14272 4372 14296 4428
rect 14352 4372 14376 4428
rect 14432 4372 14456 4428
rect 14512 4372 16740 4428
rect 11284 4368 16740 4372
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4428 28740 4432
rect 23284 4372 24216 4428
rect 24272 4372 24296 4428
rect 24352 4372 24376 4428
rect 24432 4372 24456 4428
rect 24512 4372 28740 4428
rect 23284 4368 28740 4372
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4428 34740 4432
rect 29284 4372 34216 4428
rect 34272 4372 34296 4428
rect 34352 4372 34376 4428
rect 34432 4372 34456 4428
rect 34512 4372 34740 4428
rect 29284 4368 34740 4372
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4428 46740 4432
rect 41284 4372 44216 4428
rect 44272 4372 44296 4428
rect 44352 4372 44376 4428
rect 44432 4372 44456 4428
rect 44512 4372 46740 4428
rect 41284 4368 46740 4372
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4428 58740 4432
rect 53284 4372 54216 4428
rect 54272 4372 54296 4428
rect 54352 4372 54376 4428
rect 54432 4372 54456 4428
rect 54512 4372 58740 4428
rect 53284 4368 58740 4372
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4428 64740 4432
rect 59284 4372 64216 4428
rect 64272 4372 64296 4428
rect 64352 4372 64376 4428
rect 64432 4372 64456 4428
rect 64512 4372 64740 4428
rect 59284 4368 64740 4372
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4428 75028 4432
rect 71284 4372 74216 4428
rect 74272 4372 74296 4428
rect 74352 4372 74376 4428
rect 74432 4372 74456 4428
rect 74512 4372 75028 4428
rect 71284 4368 75028 4372
rect 964 4352 75028 4368
rect 964 4348 4740 4352
rect 964 4292 4216 4348
rect 4272 4292 4296 4348
rect 4352 4292 4376 4348
rect 4432 4292 4456 4348
rect 4512 4292 4740 4348
rect 964 4288 4740 4292
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4348 16740 4352
rect 11284 4292 14216 4348
rect 14272 4292 14296 4348
rect 14352 4292 14376 4348
rect 14432 4292 14456 4348
rect 14512 4292 16740 4348
rect 11284 4288 16740 4292
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4348 28740 4352
rect 23284 4292 24216 4348
rect 24272 4292 24296 4348
rect 24352 4292 24376 4348
rect 24432 4292 24456 4348
rect 24512 4292 28740 4348
rect 23284 4288 28740 4292
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4348 34740 4352
rect 29284 4292 34216 4348
rect 34272 4292 34296 4348
rect 34352 4292 34376 4348
rect 34432 4292 34456 4348
rect 34512 4292 34740 4348
rect 29284 4288 34740 4292
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4348 46740 4352
rect 41284 4292 44216 4348
rect 44272 4292 44296 4348
rect 44352 4292 44376 4348
rect 44432 4292 44456 4348
rect 44512 4292 46740 4348
rect 41284 4288 46740 4292
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4348 58740 4352
rect 53284 4292 54216 4348
rect 54272 4292 54296 4348
rect 54352 4292 54376 4348
rect 54432 4292 54456 4348
rect 54512 4292 58740 4348
rect 53284 4288 58740 4292
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4348 64740 4352
rect 59284 4292 64216 4348
rect 64272 4292 64296 4348
rect 64352 4292 64376 4348
rect 64432 4292 64456 4348
rect 64512 4292 64740 4348
rect 59284 4288 64740 4292
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4348 75028 4352
rect 71284 4292 74216 4348
rect 74272 4292 74296 4348
rect 74352 4292 74376 4348
rect 74432 4292 74456 4348
rect 74512 4292 75028 4348
rect 71284 4288 75028 4292
rect 964 4264 75028 4288
rect 61009 4178 61075 4181
rect 61469 4178 61535 4181
rect 61009 4176 61535 4178
rect 61009 4120 61014 4176
rect 61070 4120 61474 4176
rect 61530 4120 61535 4176
rect 61009 4118 61535 4120
rect 61009 4115 61075 4118
rect 61469 4115 61535 4118
rect 31293 4042 31359 4045
rect 63718 4042 63724 4044
rect 31293 4040 63724 4042
rect 31293 3984 31298 4040
rect 31354 3984 63724 4040
rect 31293 3982 63724 3984
rect 31293 3979 31359 3982
rect 63718 3980 63724 3982
rect 63788 3980 63794 4044
rect 32765 3634 32831 3637
rect 36077 3634 36143 3637
rect 32765 3632 36143 3634
rect 32765 3576 32770 3632
rect 32826 3576 36082 3632
rect 36138 3576 36143 3632
rect 32765 3574 36143 3576
rect 32765 3571 32831 3574
rect 36077 3571 36143 3574
rect 25497 3498 25563 3501
rect 28165 3498 28231 3501
rect 25497 3496 28231 3498
rect 25497 3440 25502 3496
rect 25558 3440 28170 3496
rect 28226 3440 28231 3496
rect 25497 3438 28231 3440
rect 25497 3435 25563 3438
rect 28165 3435 28231 3438
rect 31293 3498 31359 3501
rect 33225 3498 33291 3501
rect 31293 3496 33291 3498
rect 31293 3440 31298 3496
rect 31354 3440 33230 3496
rect 33286 3440 33291 3496
rect 31293 3438 33291 3440
rect 31293 3435 31359 3438
rect 33225 3435 33291 3438
rect 14733 3362 14799 3365
rect 39982 3362 39988 3364
rect 14733 3360 39988 3362
rect 14733 3304 14738 3360
rect 14794 3304 39988 3360
rect 14733 3302 39988 3304
rect 14733 3299 14799 3302
rect 39982 3300 39988 3302
rect 40052 3300 40058 3364
rect 47853 3362 47919 3365
rect 66294 3362 66300 3364
rect 47853 3360 66300 3362
rect 47853 3304 47858 3360
rect 47914 3304 66300 3360
rect 47853 3302 66300 3304
rect 47853 3299 47919 3302
rect 66294 3300 66300 3302
rect 66364 3300 66370 3364
rect 32213 3090 32279 3093
rect 64873 3090 64939 3093
rect 32213 3088 64939 3090
rect 32213 3032 32218 3088
rect 32274 3032 64878 3088
rect 64934 3032 64939 3088
rect 32213 3030 64939 3032
rect 32213 3027 32279 3030
rect 64873 3027 64939 3030
rect 964 2240 75028 2264
rect 964 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2236 1900 2240
rect 1964 2236 1980 2240
rect 2044 2236 2060 2240
rect 2124 2236 2140 2240
rect 1884 2176 1900 2180
rect 1964 2176 1980 2180
rect 2044 2176 2060 2180
rect 2124 2176 2140 2180
rect 2204 2176 2220 2240
rect 2284 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2236 13740 2240
rect 8284 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 13740 2236
rect 8284 2176 13740 2180
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2236 25740 2240
rect 20284 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 25740 2236
rect 20284 2176 25740 2180
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2236 31900 2240
rect 31964 2236 31980 2240
rect 32044 2236 32060 2240
rect 32124 2236 32140 2240
rect 31884 2176 31900 2180
rect 31964 2176 31980 2180
rect 32044 2176 32060 2180
rect 32124 2176 32140 2180
rect 32204 2176 32220 2240
rect 32284 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2236 43740 2240
rect 38284 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 43740 2236
rect 38284 2176 43740 2180
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2236 55740 2240
rect 50284 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 55740 2236
rect 50284 2176 55740 2180
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2236 61900 2240
rect 61964 2236 61980 2240
rect 62044 2236 62060 2240
rect 62124 2236 62140 2240
rect 61884 2176 61900 2180
rect 61964 2176 61980 2180
rect 62044 2176 62060 2180
rect 62124 2176 62140 2180
rect 62204 2176 62220 2240
rect 62284 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2236 73740 2240
rect 68284 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 73740 2236
rect 68284 2176 73740 2180
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 75028 2240
rect 964 2160 75028 2176
rect 964 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2156 1900 2160
rect 1964 2156 1980 2160
rect 2044 2156 2060 2160
rect 2124 2156 2140 2160
rect 1884 2096 1900 2100
rect 1964 2096 1980 2100
rect 2044 2096 2060 2100
rect 2124 2096 2140 2100
rect 2204 2096 2220 2160
rect 2284 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2156 13740 2160
rect 8284 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 13740 2156
rect 8284 2096 13740 2100
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2156 25740 2160
rect 20284 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 25740 2156
rect 20284 2096 25740 2100
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2156 31900 2160
rect 31964 2156 31980 2160
rect 32044 2156 32060 2160
rect 32124 2156 32140 2160
rect 31884 2096 31900 2100
rect 31964 2096 31980 2100
rect 32044 2096 32060 2100
rect 32124 2096 32140 2100
rect 32204 2096 32220 2160
rect 32284 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2156 43740 2160
rect 38284 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 43740 2156
rect 38284 2096 43740 2100
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2156 55740 2160
rect 50284 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 55740 2156
rect 50284 2096 55740 2100
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2156 61900 2160
rect 61964 2156 61980 2160
rect 62044 2156 62060 2160
rect 62124 2156 62140 2160
rect 61884 2096 61900 2100
rect 61964 2096 61980 2100
rect 62044 2096 62060 2100
rect 62124 2096 62140 2100
rect 62204 2096 62220 2160
rect 62284 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2156 73740 2160
rect 68284 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 73740 2156
rect 68284 2096 73740 2100
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 75028 2160
rect 964 2080 75028 2096
rect 964 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2076 1900 2080
rect 1964 2076 1980 2080
rect 2044 2076 2060 2080
rect 2124 2076 2140 2080
rect 1884 2016 1900 2020
rect 1964 2016 1980 2020
rect 2044 2016 2060 2020
rect 2124 2016 2140 2020
rect 2204 2016 2220 2080
rect 2284 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2076 13740 2080
rect 8284 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 13740 2076
rect 8284 2016 13740 2020
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2076 25740 2080
rect 20284 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 25740 2076
rect 20284 2016 25740 2020
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2076 31900 2080
rect 31964 2076 31980 2080
rect 32044 2076 32060 2080
rect 32124 2076 32140 2080
rect 31884 2016 31900 2020
rect 31964 2016 31980 2020
rect 32044 2016 32060 2020
rect 32124 2016 32140 2020
rect 32204 2016 32220 2080
rect 32284 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2076 43740 2080
rect 38284 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 43740 2076
rect 38284 2016 43740 2020
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2076 55740 2080
rect 50284 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 55740 2076
rect 50284 2016 55740 2020
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2076 61900 2080
rect 61964 2076 61980 2080
rect 62044 2076 62060 2080
rect 62124 2076 62140 2080
rect 61884 2016 61900 2020
rect 61964 2016 61980 2020
rect 62044 2016 62060 2020
rect 62124 2016 62140 2020
rect 62204 2016 62220 2080
rect 62284 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2076 73740 2080
rect 68284 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 73740 2076
rect 68284 2016 73740 2020
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 75028 2080
rect 964 2000 75028 2016
rect 964 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1996 1900 2000
rect 1964 1996 1980 2000
rect 2044 1996 2060 2000
rect 2124 1996 2140 2000
rect 1884 1936 1900 1940
rect 1964 1936 1980 1940
rect 2044 1936 2060 1940
rect 2124 1936 2140 1940
rect 2204 1936 2220 2000
rect 2284 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1996 13740 2000
rect 8284 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 13740 1996
rect 8284 1936 13740 1940
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1996 25740 2000
rect 20284 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 25740 1996
rect 20284 1936 25740 1940
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1996 31900 2000
rect 31964 1996 31980 2000
rect 32044 1996 32060 2000
rect 32124 1996 32140 2000
rect 31884 1936 31900 1940
rect 31964 1936 31980 1940
rect 32044 1936 32060 1940
rect 32124 1936 32140 1940
rect 32204 1936 32220 2000
rect 32284 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1996 43740 2000
rect 38284 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 43740 1996
rect 38284 1936 43740 1940
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1996 55740 2000
rect 50284 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 55740 1996
rect 50284 1936 55740 1940
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1996 61900 2000
rect 61964 1996 61980 2000
rect 62044 1996 62060 2000
rect 62124 1996 62140 2000
rect 61884 1936 61900 1940
rect 61964 1936 61980 1940
rect 62044 1936 62060 1940
rect 62124 1936 62140 1940
rect 62204 1936 62220 2000
rect 62284 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1996 73740 2000
rect 68284 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 73740 1996
rect 68284 1936 73740 1940
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 75028 2000
rect 964 1912 75028 1936
<< via3 >>
rect 4740 84528 4804 84592
rect 4820 84528 4884 84592
rect 4900 84528 4964 84592
rect 4980 84528 5044 84592
rect 5060 84528 5124 84592
rect 5140 84528 5204 84592
rect 5220 84528 5284 84592
rect 10740 84528 10804 84592
rect 10820 84528 10884 84592
rect 10900 84528 10964 84592
rect 10980 84528 11044 84592
rect 11060 84528 11124 84592
rect 11140 84528 11204 84592
rect 11220 84528 11284 84592
rect 16740 84528 16804 84592
rect 16820 84528 16884 84592
rect 16900 84528 16964 84592
rect 16980 84528 17044 84592
rect 17060 84528 17124 84592
rect 17140 84528 17204 84592
rect 17220 84528 17284 84592
rect 22740 84528 22804 84592
rect 22820 84528 22884 84592
rect 22900 84528 22964 84592
rect 22980 84528 23044 84592
rect 23060 84528 23124 84592
rect 23140 84528 23204 84592
rect 23220 84528 23284 84592
rect 28740 84528 28804 84592
rect 28820 84528 28884 84592
rect 28900 84528 28964 84592
rect 28980 84528 29044 84592
rect 29060 84528 29124 84592
rect 29140 84528 29204 84592
rect 29220 84528 29284 84592
rect 34740 84528 34804 84592
rect 34820 84528 34884 84592
rect 34900 84528 34964 84592
rect 34980 84528 35044 84592
rect 35060 84528 35124 84592
rect 35140 84528 35204 84592
rect 35220 84528 35284 84592
rect 40740 84528 40804 84592
rect 40820 84528 40884 84592
rect 40900 84528 40964 84592
rect 40980 84528 41044 84592
rect 41060 84528 41124 84592
rect 41140 84528 41204 84592
rect 41220 84528 41284 84592
rect 46740 84528 46804 84592
rect 46820 84528 46884 84592
rect 46900 84528 46964 84592
rect 46980 84528 47044 84592
rect 47060 84528 47124 84592
rect 47140 84528 47204 84592
rect 47220 84528 47284 84592
rect 52740 84528 52804 84592
rect 52820 84528 52884 84592
rect 52900 84528 52964 84592
rect 52980 84528 53044 84592
rect 53060 84528 53124 84592
rect 53140 84528 53204 84592
rect 53220 84528 53284 84592
rect 58740 84528 58804 84592
rect 58820 84528 58884 84592
rect 58900 84528 58964 84592
rect 58980 84528 59044 84592
rect 59060 84528 59124 84592
rect 59140 84528 59204 84592
rect 59220 84528 59284 84592
rect 64740 84528 64804 84592
rect 64820 84528 64884 84592
rect 64900 84528 64964 84592
rect 64980 84528 65044 84592
rect 65060 84528 65124 84592
rect 65140 84528 65204 84592
rect 65220 84528 65284 84592
rect 70740 84528 70804 84592
rect 70820 84528 70884 84592
rect 70900 84528 70964 84592
rect 70980 84528 71044 84592
rect 71060 84528 71124 84592
rect 71140 84528 71204 84592
rect 71220 84528 71284 84592
rect 4740 84448 4804 84512
rect 4820 84448 4884 84512
rect 4900 84448 4964 84512
rect 4980 84448 5044 84512
rect 5060 84448 5124 84512
rect 5140 84448 5204 84512
rect 5220 84448 5284 84512
rect 10740 84448 10804 84512
rect 10820 84448 10884 84512
rect 10900 84448 10964 84512
rect 10980 84448 11044 84512
rect 11060 84448 11124 84512
rect 11140 84448 11204 84512
rect 11220 84448 11284 84512
rect 16740 84448 16804 84512
rect 16820 84448 16884 84512
rect 16900 84448 16964 84512
rect 16980 84448 17044 84512
rect 17060 84448 17124 84512
rect 17140 84448 17204 84512
rect 17220 84448 17284 84512
rect 22740 84448 22804 84512
rect 22820 84448 22884 84512
rect 22900 84448 22964 84512
rect 22980 84448 23044 84512
rect 23060 84448 23124 84512
rect 23140 84448 23204 84512
rect 23220 84448 23284 84512
rect 28740 84448 28804 84512
rect 28820 84448 28884 84512
rect 28900 84448 28964 84512
rect 28980 84448 29044 84512
rect 29060 84448 29124 84512
rect 29140 84448 29204 84512
rect 29220 84448 29284 84512
rect 34740 84448 34804 84512
rect 34820 84448 34884 84512
rect 34900 84448 34964 84512
rect 34980 84448 35044 84512
rect 35060 84448 35124 84512
rect 35140 84448 35204 84512
rect 35220 84448 35284 84512
rect 40740 84448 40804 84512
rect 40820 84448 40884 84512
rect 40900 84448 40964 84512
rect 40980 84448 41044 84512
rect 41060 84448 41124 84512
rect 41140 84448 41204 84512
rect 41220 84448 41284 84512
rect 46740 84448 46804 84512
rect 46820 84448 46884 84512
rect 46900 84448 46964 84512
rect 46980 84448 47044 84512
rect 47060 84448 47124 84512
rect 47140 84448 47204 84512
rect 47220 84448 47284 84512
rect 52740 84448 52804 84512
rect 52820 84448 52884 84512
rect 52900 84448 52964 84512
rect 52980 84448 53044 84512
rect 53060 84448 53124 84512
rect 53140 84448 53204 84512
rect 53220 84448 53284 84512
rect 58740 84448 58804 84512
rect 58820 84448 58884 84512
rect 58900 84448 58964 84512
rect 58980 84448 59044 84512
rect 59060 84448 59124 84512
rect 59140 84448 59204 84512
rect 59220 84448 59284 84512
rect 64740 84448 64804 84512
rect 64820 84448 64884 84512
rect 64900 84448 64964 84512
rect 64980 84448 65044 84512
rect 65060 84448 65124 84512
rect 65140 84448 65204 84512
rect 65220 84448 65284 84512
rect 70740 84448 70804 84512
rect 70820 84448 70884 84512
rect 70900 84448 70964 84512
rect 70980 84448 71044 84512
rect 71060 84448 71124 84512
rect 71140 84448 71204 84512
rect 71220 84448 71284 84512
rect 4740 84368 4804 84432
rect 4820 84368 4884 84432
rect 4900 84368 4964 84432
rect 4980 84368 5044 84432
rect 5060 84368 5124 84432
rect 5140 84368 5204 84432
rect 5220 84368 5284 84432
rect 10740 84368 10804 84432
rect 10820 84368 10884 84432
rect 10900 84368 10964 84432
rect 10980 84368 11044 84432
rect 11060 84368 11124 84432
rect 11140 84368 11204 84432
rect 11220 84368 11284 84432
rect 16740 84368 16804 84432
rect 16820 84368 16884 84432
rect 16900 84368 16964 84432
rect 16980 84368 17044 84432
rect 17060 84368 17124 84432
rect 17140 84368 17204 84432
rect 17220 84368 17284 84432
rect 22740 84368 22804 84432
rect 22820 84368 22884 84432
rect 22900 84368 22964 84432
rect 22980 84368 23044 84432
rect 23060 84368 23124 84432
rect 23140 84368 23204 84432
rect 23220 84368 23284 84432
rect 28740 84368 28804 84432
rect 28820 84368 28884 84432
rect 28900 84368 28964 84432
rect 28980 84368 29044 84432
rect 29060 84368 29124 84432
rect 29140 84368 29204 84432
rect 29220 84368 29284 84432
rect 34740 84368 34804 84432
rect 34820 84368 34884 84432
rect 34900 84368 34964 84432
rect 34980 84368 35044 84432
rect 35060 84368 35124 84432
rect 35140 84368 35204 84432
rect 35220 84368 35284 84432
rect 40740 84368 40804 84432
rect 40820 84368 40884 84432
rect 40900 84368 40964 84432
rect 40980 84368 41044 84432
rect 41060 84368 41124 84432
rect 41140 84368 41204 84432
rect 41220 84368 41284 84432
rect 46740 84368 46804 84432
rect 46820 84368 46884 84432
rect 46900 84368 46964 84432
rect 46980 84368 47044 84432
rect 47060 84368 47124 84432
rect 47140 84368 47204 84432
rect 47220 84368 47284 84432
rect 52740 84368 52804 84432
rect 52820 84368 52884 84432
rect 52900 84368 52964 84432
rect 52980 84368 53044 84432
rect 53060 84368 53124 84432
rect 53140 84368 53204 84432
rect 53220 84368 53284 84432
rect 58740 84368 58804 84432
rect 58820 84368 58884 84432
rect 58900 84368 58964 84432
rect 58980 84368 59044 84432
rect 59060 84368 59124 84432
rect 59140 84368 59204 84432
rect 59220 84368 59284 84432
rect 64740 84368 64804 84432
rect 64820 84368 64884 84432
rect 64900 84368 64964 84432
rect 64980 84368 65044 84432
rect 65060 84368 65124 84432
rect 65140 84368 65204 84432
rect 65220 84368 65284 84432
rect 70740 84368 70804 84432
rect 70820 84368 70884 84432
rect 70900 84368 70964 84432
rect 70980 84368 71044 84432
rect 71060 84368 71124 84432
rect 71140 84368 71204 84432
rect 71220 84368 71284 84432
rect 4740 84288 4804 84352
rect 4820 84288 4884 84352
rect 4900 84288 4964 84352
rect 4980 84288 5044 84352
rect 5060 84288 5124 84352
rect 5140 84288 5204 84352
rect 5220 84288 5284 84352
rect 10740 84288 10804 84352
rect 10820 84288 10884 84352
rect 10900 84288 10964 84352
rect 10980 84288 11044 84352
rect 11060 84288 11124 84352
rect 11140 84288 11204 84352
rect 11220 84288 11284 84352
rect 16740 84288 16804 84352
rect 16820 84288 16884 84352
rect 16900 84288 16964 84352
rect 16980 84288 17044 84352
rect 17060 84288 17124 84352
rect 17140 84288 17204 84352
rect 17220 84288 17284 84352
rect 22740 84288 22804 84352
rect 22820 84288 22884 84352
rect 22900 84288 22964 84352
rect 22980 84288 23044 84352
rect 23060 84288 23124 84352
rect 23140 84288 23204 84352
rect 23220 84288 23284 84352
rect 28740 84288 28804 84352
rect 28820 84288 28884 84352
rect 28900 84288 28964 84352
rect 28980 84288 29044 84352
rect 29060 84288 29124 84352
rect 29140 84288 29204 84352
rect 29220 84288 29284 84352
rect 34740 84288 34804 84352
rect 34820 84288 34884 84352
rect 34900 84288 34964 84352
rect 34980 84288 35044 84352
rect 35060 84288 35124 84352
rect 35140 84288 35204 84352
rect 35220 84288 35284 84352
rect 40740 84288 40804 84352
rect 40820 84288 40884 84352
rect 40900 84288 40964 84352
rect 40980 84288 41044 84352
rect 41060 84288 41124 84352
rect 41140 84288 41204 84352
rect 41220 84288 41284 84352
rect 46740 84288 46804 84352
rect 46820 84288 46884 84352
rect 46900 84288 46964 84352
rect 46980 84288 47044 84352
rect 47060 84288 47124 84352
rect 47140 84288 47204 84352
rect 47220 84288 47284 84352
rect 52740 84288 52804 84352
rect 52820 84288 52884 84352
rect 52900 84288 52964 84352
rect 52980 84288 53044 84352
rect 53060 84288 53124 84352
rect 53140 84288 53204 84352
rect 53220 84288 53284 84352
rect 58740 84288 58804 84352
rect 58820 84288 58884 84352
rect 58900 84288 58964 84352
rect 58980 84288 59044 84352
rect 59060 84288 59124 84352
rect 59140 84288 59204 84352
rect 59220 84288 59284 84352
rect 64740 84288 64804 84352
rect 64820 84288 64884 84352
rect 64900 84288 64964 84352
rect 64980 84288 65044 84352
rect 65060 84288 65124 84352
rect 65140 84288 65204 84352
rect 65220 84288 65284 84352
rect 70740 84288 70804 84352
rect 70820 84288 70884 84352
rect 70900 84288 70964 84352
rect 70980 84288 71044 84352
rect 71060 84288 71124 84352
rect 71140 84288 71204 84352
rect 71220 84288 71284 84352
rect 1740 82176 1804 82240
rect 1820 82176 1884 82240
rect 1900 82176 1964 82240
rect 1980 82176 2044 82240
rect 2060 82176 2124 82240
rect 2140 82176 2204 82240
rect 2220 82176 2284 82240
rect 7740 82176 7804 82240
rect 7820 82176 7884 82240
rect 7900 82176 7964 82240
rect 7980 82176 8044 82240
rect 8060 82176 8124 82240
rect 8140 82176 8204 82240
rect 8220 82176 8284 82240
rect 13740 82176 13804 82240
rect 13820 82176 13884 82240
rect 13900 82176 13964 82240
rect 13980 82176 14044 82240
rect 14060 82176 14124 82240
rect 14140 82176 14204 82240
rect 14220 82176 14284 82240
rect 19740 82176 19804 82240
rect 19820 82176 19884 82240
rect 19900 82176 19964 82240
rect 19980 82176 20044 82240
rect 20060 82176 20124 82240
rect 20140 82176 20204 82240
rect 20220 82176 20284 82240
rect 25740 82176 25804 82240
rect 25820 82176 25884 82240
rect 25900 82176 25964 82240
rect 25980 82176 26044 82240
rect 26060 82176 26124 82240
rect 26140 82176 26204 82240
rect 26220 82176 26284 82240
rect 31740 82176 31804 82240
rect 31820 82176 31884 82240
rect 31900 82176 31964 82240
rect 31980 82176 32044 82240
rect 32060 82176 32124 82240
rect 32140 82176 32204 82240
rect 32220 82176 32284 82240
rect 37740 82176 37804 82240
rect 37820 82176 37884 82240
rect 37900 82176 37964 82240
rect 37980 82176 38044 82240
rect 38060 82176 38124 82240
rect 38140 82176 38204 82240
rect 38220 82176 38284 82240
rect 43740 82176 43804 82240
rect 43820 82176 43884 82240
rect 43900 82176 43964 82240
rect 43980 82176 44044 82240
rect 44060 82176 44124 82240
rect 44140 82176 44204 82240
rect 44220 82176 44284 82240
rect 49740 82176 49804 82240
rect 49820 82176 49884 82240
rect 49900 82176 49964 82240
rect 49980 82176 50044 82240
rect 50060 82176 50124 82240
rect 50140 82176 50204 82240
rect 50220 82176 50284 82240
rect 55740 82176 55804 82240
rect 55820 82176 55884 82240
rect 55900 82176 55964 82240
rect 55980 82176 56044 82240
rect 56060 82176 56124 82240
rect 56140 82176 56204 82240
rect 56220 82176 56284 82240
rect 61740 82176 61804 82240
rect 61820 82176 61884 82240
rect 61900 82176 61964 82240
rect 61980 82176 62044 82240
rect 62060 82176 62124 82240
rect 62140 82176 62204 82240
rect 62220 82176 62284 82240
rect 67740 82176 67804 82240
rect 67820 82176 67884 82240
rect 67900 82176 67964 82240
rect 67980 82176 68044 82240
rect 68060 82176 68124 82240
rect 68140 82176 68204 82240
rect 68220 82176 68284 82240
rect 73740 82176 73804 82240
rect 73820 82176 73884 82240
rect 73900 82176 73964 82240
rect 73980 82176 74044 82240
rect 74060 82176 74124 82240
rect 74140 82176 74204 82240
rect 74220 82176 74284 82240
rect 1740 82096 1804 82160
rect 1820 82096 1884 82160
rect 1900 82096 1964 82160
rect 1980 82096 2044 82160
rect 2060 82096 2124 82160
rect 2140 82096 2204 82160
rect 2220 82096 2284 82160
rect 7740 82096 7804 82160
rect 7820 82096 7884 82160
rect 7900 82096 7964 82160
rect 7980 82096 8044 82160
rect 8060 82096 8124 82160
rect 8140 82096 8204 82160
rect 8220 82096 8284 82160
rect 13740 82096 13804 82160
rect 13820 82096 13884 82160
rect 13900 82096 13964 82160
rect 13980 82096 14044 82160
rect 14060 82096 14124 82160
rect 14140 82096 14204 82160
rect 14220 82096 14284 82160
rect 19740 82096 19804 82160
rect 19820 82096 19884 82160
rect 19900 82096 19964 82160
rect 19980 82096 20044 82160
rect 20060 82096 20124 82160
rect 20140 82096 20204 82160
rect 20220 82096 20284 82160
rect 25740 82096 25804 82160
rect 25820 82096 25884 82160
rect 25900 82096 25964 82160
rect 25980 82096 26044 82160
rect 26060 82096 26124 82160
rect 26140 82096 26204 82160
rect 26220 82096 26284 82160
rect 31740 82096 31804 82160
rect 31820 82096 31884 82160
rect 31900 82096 31964 82160
rect 31980 82096 32044 82160
rect 32060 82096 32124 82160
rect 32140 82096 32204 82160
rect 32220 82096 32284 82160
rect 37740 82096 37804 82160
rect 37820 82096 37884 82160
rect 37900 82096 37964 82160
rect 37980 82096 38044 82160
rect 38060 82096 38124 82160
rect 38140 82096 38204 82160
rect 38220 82096 38284 82160
rect 43740 82096 43804 82160
rect 43820 82096 43884 82160
rect 43900 82096 43964 82160
rect 43980 82096 44044 82160
rect 44060 82096 44124 82160
rect 44140 82096 44204 82160
rect 44220 82096 44284 82160
rect 49740 82096 49804 82160
rect 49820 82096 49884 82160
rect 49900 82096 49964 82160
rect 49980 82096 50044 82160
rect 50060 82096 50124 82160
rect 50140 82096 50204 82160
rect 50220 82096 50284 82160
rect 55740 82096 55804 82160
rect 55820 82096 55884 82160
rect 55900 82096 55964 82160
rect 55980 82096 56044 82160
rect 56060 82096 56124 82160
rect 56140 82096 56204 82160
rect 56220 82096 56284 82160
rect 61740 82096 61804 82160
rect 61820 82096 61884 82160
rect 61900 82096 61964 82160
rect 61980 82096 62044 82160
rect 62060 82096 62124 82160
rect 62140 82096 62204 82160
rect 62220 82096 62284 82160
rect 67740 82096 67804 82160
rect 67820 82096 67884 82160
rect 67900 82096 67964 82160
rect 67980 82096 68044 82160
rect 68060 82096 68124 82160
rect 68140 82096 68204 82160
rect 68220 82096 68284 82160
rect 73740 82096 73804 82160
rect 73820 82096 73884 82160
rect 73900 82096 73964 82160
rect 73980 82096 74044 82160
rect 74060 82096 74124 82160
rect 74140 82096 74204 82160
rect 74220 82096 74284 82160
rect 1740 82016 1804 82080
rect 1820 82016 1884 82080
rect 1900 82016 1964 82080
rect 1980 82016 2044 82080
rect 2060 82016 2124 82080
rect 2140 82016 2204 82080
rect 2220 82016 2284 82080
rect 7740 82016 7804 82080
rect 7820 82016 7884 82080
rect 7900 82016 7964 82080
rect 7980 82016 8044 82080
rect 8060 82016 8124 82080
rect 8140 82016 8204 82080
rect 8220 82016 8284 82080
rect 13740 82016 13804 82080
rect 13820 82016 13884 82080
rect 13900 82016 13964 82080
rect 13980 82016 14044 82080
rect 14060 82016 14124 82080
rect 14140 82016 14204 82080
rect 14220 82016 14284 82080
rect 19740 82016 19804 82080
rect 19820 82016 19884 82080
rect 19900 82016 19964 82080
rect 19980 82016 20044 82080
rect 20060 82016 20124 82080
rect 20140 82016 20204 82080
rect 20220 82016 20284 82080
rect 25740 82016 25804 82080
rect 25820 82016 25884 82080
rect 25900 82016 25964 82080
rect 25980 82016 26044 82080
rect 26060 82016 26124 82080
rect 26140 82016 26204 82080
rect 26220 82016 26284 82080
rect 31740 82016 31804 82080
rect 31820 82016 31884 82080
rect 31900 82016 31964 82080
rect 31980 82016 32044 82080
rect 32060 82016 32124 82080
rect 32140 82016 32204 82080
rect 32220 82016 32284 82080
rect 37740 82016 37804 82080
rect 37820 82016 37884 82080
rect 37900 82016 37964 82080
rect 37980 82016 38044 82080
rect 38060 82016 38124 82080
rect 38140 82016 38204 82080
rect 38220 82016 38284 82080
rect 43740 82016 43804 82080
rect 43820 82016 43884 82080
rect 43900 82016 43964 82080
rect 43980 82016 44044 82080
rect 44060 82016 44124 82080
rect 44140 82016 44204 82080
rect 44220 82016 44284 82080
rect 49740 82016 49804 82080
rect 49820 82016 49884 82080
rect 49900 82016 49964 82080
rect 49980 82016 50044 82080
rect 50060 82016 50124 82080
rect 50140 82016 50204 82080
rect 50220 82016 50284 82080
rect 55740 82016 55804 82080
rect 55820 82016 55884 82080
rect 55900 82016 55964 82080
rect 55980 82016 56044 82080
rect 56060 82016 56124 82080
rect 56140 82016 56204 82080
rect 56220 82016 56284 82080
rect 61740 82016 61804 82080
rect 61820 82016 61884 82080
rect 61900 82016 61964 82080
rect 61980 82016 62044 82080
rect 62060 82016 62124 82080
rect 62140 82016 62204 82080
rect 62220 82016 62284 82080
rect 67740 82016 67804 82080
rect 67820 82016 67884 82080
rect 67900 82016 67964 82080
rect 67980 82016 68044 82080
rect 68060 82016 68124 82080
rect 68140 82016 68204 82080
rect 68220 82016 68284 82080
rect 73740 82016 73804 82080
rect 73820 82016 73884 82080
rect 73900 82016 73964 82080
rect 73980 82016 74044 82080
rect 74060 82016 74124 82080
rect 74140 82016 74204 82080
rect 74220 82016 74284 82080
rect 1740 81936 1804 82000
rect 1820 81936 1884 82000
rect 1900 81936 1964 82000
rect 1980 81936 2044 82000
rect 2060 81936 2124 82000
rect 2140 81936 2204 82000
rect 2220 81936 2284 82000
rect 7740 81936 7804 82000
rect 7820 81936 7884 82000
rect 7900 81936 7964 82000
rect 7980 81936 8044 82000
rect 8060 81936 8124 82000
rect 8140 81936 8204 82000
rect 8220 81936 8284 82000
rect 13740 81936 13804 82000
rect 13820 81936 13884 82000
rect 13900 81936 13964 82000
rect 13980 81936 14044 82000
rect 14060 81936 14124 82000
rect 14140 81936 14204 82000
rect 14220 81936 14284 82000
rect 19740 81936 19804 82000
rect 19820 81936 19884 82000
rect 19900 81936 19964 82000
rect 19980 81936 20044 82000
rect 20060 81936 20124 82000
rect 20140 81936 20204 82000
rect 20220 81936 20284 82000
rect 25740 81936 25804 82000
rect 25820 81936 25884 82000
rect 25900 81936 25964 82000
rect 25980 81936 26044 82000
rect 26060 81936 26124 82000
rect 26140 81936 26204 82000
rect 26220 81936 26284 82000
rect 31740 81936 31804 82000
rect 31820 81936 31884 82000
rect 31900 81936 31964 82000
rect 31980 81936 32044 82000
rect 32060 81936 32124 82000
rect 32140 81936 32204 82000
rect 32220 81936 32284 82000
rect 37740 81936 37804 82000
rect 37820 81936 37884 82000
rect 37900 81936 37964 82000
rect 37980 81936 38044 82000
rect 38060 81936 38124 82000
rect 38140 81936 38204 82000
rect 38220 81936 38284 82000
rect 43740 81936 43804 82000
rect 43820 81936 43884 82000
rect 43900 81936 43964 82000
rect 43980 81936 44044 82000
rect 44060 81936 44124 82000
rect 44140 81936 44204 82000
rect 44220 81936 44284 82000
rect 49740 81936 49804 82000
rect 49820 81936 49884 82000
rect 49900 81936 49964 82000
rect 49980 81936 50044 82000
rect 50060 81936 50124 82000
rect 50140 81936 50204 82000
rect 50220 81936 50284 82000
rect 55740 81936 55804 82000
rect 55820 81936 55884 82000
rect 55900 81936 55964 82000
rect 55980 81936 56044 82000
rect 56060 81936 56124 82000
rect 56140 81936 56204 82000
rect 56220 81936 56284 82000
rect 61740 81936 61804 82000
rect 61820 81936 61884 82000
rect 61900 81936 61964 82000
rect 61980 81936 62044 82000
rect 62060 81936 62124 82000
rect 62140 81936 62204 82000
rect 62220 81936 62284 82000
rect 67740 81936 67804 82000
rect 67820 81936 67884 82000
rect 67900 81936 67964 82000
rect 67980 81936 68044 82000
rect 68060 81936 68124 82000
rect 68140 81936 68204 82000
rect 68220 81936 68284 82000
rect 73740 81936 73804 82000
rect 73820 81936 73884 82000
rect 73900 81936 73964 82000
rect 73980 81936 74044 82000
rect 74060 81936 74124 82000
rect 74140 81936 74204 82000
rect 74220 81936 74284 82000
rect 4740 74528 4804 74592
rect 4820 74528 4884 74592
rect 4900 74528 4964 74592
rect 4980 74528 5044 74592
rect 5060 74528 5124 74592
rect 5140 74528 5204 74592
rect 5220 74528 5284 74592
rect 10740 74528 10804 74592
rect 10820 74528 10884 74592
rect 10900 74528 10964 74592
rect 10980 74528 11044 74592
rect 11060 74528 11124 74592
rect 11140 74528 11204 74592
rect 11220 74528 11284 74592
rect 16740 74528 16804 74592
rect 16820 74528 16884 74592
rect 16900 74528 16964 74592
rect 16980 74528 17044 74592
rect 17060 74528 17124 74592
rect 17140 74528 17204 74592
rect 17220 74528 17284 74592
rect 22740 74528 22804 74592
rect 22820 74528 22884 74592
rect 22900 74528 22964 74592
rect 22980 74528 23044 74592
rect 23060 74528 23124 74592
rect 23140 74528 23204 74592
rect 23220 74528 23284 74592
rect 28740 74528 28804 74592
rect 28820 74528 28884 74592
rect 28900 74528 28964 74592
rect 28980 74528 29044 74592
rect 29060 74528 29124 74592
rect 29140 74528 29204 74592
rect 29220 74528 29284 74592
rect 34740 74528 34804 74592
rect 34820 74528 34884 74592
rect 34900 74528 34964 74592
rect 34980 74528 35044 74592
rect 35060 74528 35124 74592
rect 35140 74528 35204 74592
rect 35220 74528 35284 74592
rect 40740 74528 40804 74592
rect 40820 74528 40884 74592
rect 40900 74528 40964 74592
rect 40980 74528 41044 74592
rect 41060 74528 41124 74592
rect 41140 74528 41204 74592
rect 41220 74528 41284 74592
rect 46740 74528 46804 74592
rect 46820 74528 46884 74592
rect 46900 74528 46964 74592
rect 46980 74528 47044 74592
rect 47060 74528 47124 74592
rect 47140 74528 47204 74592
rect 47220 74528 47284 74592
rect 52740 74528 52804 74592
rect 52820 74528 52884 74592
rect 52900 74528 52964 74592
rect 52980 74528 53044 74592
rect 53060 74528 53124 74592
rect 53140 74528 53204 74592
rect 53220 74528 53284 74592
rect 58740 74528 58804 74592
rect 58820 74528 58884 74592
rect 58900 74528 58964 74592
rect 58980 74528 59044 74592
rect 59060 74528 59124 74592
rect 59140 74528 59204 74592
rect 59220 74528 59284 74592
rect 64740 74528 64804 74592
rect 64820 74528 64884 74592
rect 64900 74528 64964 74592
rect 64980 74528 65044 74592
rect 65060 74528 65124 74592
rect 65140 74528 65204 74592
rect 65220 74528 65284 74592
rect 70740 74528 70804 74592
rect 70820 74528 70884 74592
rect 70900 74528 70964 74592
rect 70980 74528 71044 74592
rect 71060 74528 71124 74592
rect 71140 74528 71204 74592
rect 71220 74528 71284 74592
rect 4740 74448 4804 74512
rect 4820 74448 4884 74512
rect 4900 74448 4964 74512
rect 4980 74448 5044 74512
rect 5060 74448 5124 74512
rect 5140 74448 5204 74512
rect 5220 74448 5284 74512
rect 10740 74448 10804 74512
rect 10820 74448 10884 74512
rect 10900 74448 10964 74512
rect 10980 74448 11044 74512
rect 11060 74448 11124 74512
rect 11140 74448 11204 74512
rect 11220 74448 11284 74512
rect 16740 74448 16804 74512
rect 16820 74448 16884 74512
rect 16900 74448 16964 74512
rect 16980 74448 17044 74512
rect 17060 74448 17124 74512
rect 17140 74448 17204 74512
rect 17220 74448 17284 74512
rect 22740 74448 22804 74512
rect 22820 74448 22884 74512
rect 22900 74448 22964 74512
rect 22980 74448 23044 74512
rect 23060 74448 23124 74512
rect 23140 74448 23204 74512
rect 23220 74448 23284 74512
rect 28740 74448 28804 74512
rect 28820 74448 28884 74512
rect 28900 74448 28964 74512
rect 28980 74448 29044 74512
rect 29060 74448 29124 74512
rect 29140 74448 29204 74512
rect 29220 74448 29284 74512
rect 34740 74448 34804 74512
rect 34820 74448 34884 74512
rect 34900 74448 34964 74512
rect 34980 74448 35044 74512
rect 35060 74448 35124 74512
rect 35140 74448 35204 74512
rect 35220 74448 35284 74512
rect 40740 74448 40804 74512
rect 40820 74448 40884 74512
rect 40900 74448 40964 74512
rect 40980 74448 41044 74512
rect 41060 74448 41124 74512
rect 41140 74448 41204 74512
rect 41220 74448 41284 74512
rect 46740 74448 46804 74512
rect 46820 74448 46884 74512
rect 46900 74448 46964 74512
rect 46980 74448 47044 74512
rect 47060 74448 47124 74512
rect 47140 74448 47204 74512
rect 47220 74448 47284 74512
rect 52740 74448 52804 74512
rect 52820 74448 52884 74512
rect 52900 74448 52964 74512
rect 52980 74448 53044 74512
rect 53060 74448 53124 74512
rect 53140 74448 53204 74512
rect 53220 74448 53284 74512
rect 58740 74448 58804 74512
rect 58820 74448 58884 74512
rect 58900 74448 58964 74512
rect 58980 74448 59044 74512
rect 59060 74448 59124 74512
rect 59140 74448 59204 74512
rect 59220 74448 59284 74512
rect 64740 74448 64804 74512
rect 64820 74448 64884 74512
rect 64900 74448 64964 74512
rect 64980 74448 65044 74512
rect 65060 74448 65124 74512
rect 65140 74448 65204 74512
rect 65220 74448 65284 74512
rect 70740 74448 70804 74512
rect 70820 74448 70884 74512
rect 70900 74448 70964 74512
rect 70980 74448 71044 74512
rect 71060 74448 71124 74512
rect 71140 74448 71204 74512
rect 71220 74448 71284 74512
rect 4740 74368 4804 74432
rect 4820 74368 4884 74432
rect 4900 74368 4964 74432
rect 4980 74368 5044 74432
rect 5060 74368 5124 74432
rect 5140 74368 5204 74432
rect 5220 74368 5284 74432
rect 10740 74368 10804 74432
rect 10820 74368 10884 74432
rect 10900 74368 10964 74432
rect 10980 74368 11044 74432
rect 11060 74368 11124 74432
rect 11140 74368 11204 74432
rect 11220 74368 11284 74432
rect 16740 74368 16804 74432
rect 16820 74368 16884 74432
rect 16900 74368 16964 74432
rect 16980 74368 17044 74432
rect 17060 74368 17124 74432
rect 17140 74368 17204 74432
rect 17220 74368 17284 74432
rect 22740 74368 22804 74432
rect 22820 74368 22884 74432
rect 22900 74368 22964 74432
rect 22980 74368 23044 74432
rect 23060 74368 23124 74432
rect 23140 74368 23204 74432
rect 23220 74368 23284 74432
rect 28740 74368 28804 74432
rect 28820 74368 28884 74432
rect 28900 74368 28964 74432
rect 28980 74368 29044 74432
rect 29060 74368 29124 74432
rect 29140 74368 29204 74432
rect 29220 74368 29284 74432
rect 34740 74368 34804 74432
rect 34820 74368 34884 74432
rect 34900 74368 34964 74432
rect 34980 74368 35044 74432
rect 35060 74368 35124 74432
rect 35140 74368 35204 74432
rect 35220 74368 35284 74432
rect 40740 74368 40804 74432
rect 40820 74368 40884 74432
rect 40900 74368 40964 74432
rect 40980 74368 41044 74432
rect 41060 74368 41124 74432
rect 41140 74368 41204 74432
rect 41220 74368 41284 74432
rect 46740 74368 46804 74432
rect 46820 74368 46884 74432
rect 46900 74368 46964 74432
rect 46980 74368 47044 74432
rect 47060 74368 47124 74432
rect 47140 74368 47204 74432
rect 47220 74368 47284 74432
rect 52740 74368 52804 74432
rect 52820 74368 52884 74432
rect 52900 74368 52964 74432
rect 52980 74368 53044 74432
rect 53060 74368 53124 74432
rect 53140 74368 53204 74432
rect 53220 74368 53284 74432
rect 58740 74368 58804 74432
rect 58820 74368 58884 74432
rect 58900 74368 58964 74432
rect 58980 74368 59044 74432
rect 59060 74368 59124 74432
rect 59140 74368 59204 74432
rect 59220 74368 59284 74432
rect 64740 74368 64804 74432
rect 64820 74368 64884 74432
rect 64900 74368 64964 74432
rect 64980 74368 65044 74432
rect 65060 74368 65124 74432
rect 65140 74368 65204 74432
rect 65220 74368 65284 74432
rect 70740 74368 70804 74432
rect 70820 74368 70884 74432
rect 70900 74368 70964 74432
rect 70980 74368 71044 74432
rect 71060 74368 71124 74432
rect 71140 74368 71204 74432
rect 71220 74368 71284 74432
rect 4740 74288 4804 74352
rect 4820 74288 4884 74352
rect 4900 74288 4964 74352
rect 4980 74288 5044 74352
rect 5060 74288 5124 74352
rect 5140 74288 5204 74352
rect 5220 74288 5284 74352
rect 10740 74288 10804 74352
rect 10820 74288 10884 74352
rect 10900 74288 10964 74352
rect 10980 74288 11044 74352
rect 11060 74288 11124 74352
rect 11140 74288 11204 74352
rect 11220 74288 11284 74352
rect 16740 74288 16804 74352
rect 16820 74288 16884 74352
rect 16900 74288 16964 74352
rect 16980 74288 17044 74352
rect 17060 74288 17124 74352
rect 17140 74288 17204 74352
rect 17220 74288 17284 74352
rect 22740 74288 22804 74352
rect 22820 74288 22884 74352
rect 22900 74288 22964 74352
rect 22980 74288 23044 74352
rect 23060 74288 23124 74352
rect 23140 74288 23204 74352
rect 23220 74288 23284 74352
rect 28740 74288 28804 74352
rect 28820 74288 28884 74352
rect 28900 74288 28964 74352
rect 28980 74288 29044 74352
rect 29060 74288 29124 74352
rect 29140 74288 29204 74352
rect 29220 74288 29284 74352
rect 34740 74288 34804 74352
rect 34820 74288 34884 74352
rect 34900 74288 34964 74352
rect 34980 74288 35044 74352
rect 35060 74288 35124 74352
rect 35140 74288 35204 74352
rect 35220 74288 35284 74352
rect 40740 74288 40804 74352
rect 40820 74288 40884 74352
rect 40900 74288 40964 74352
rect 40980 74288 41044 74352
rect 41060 74288 41124 74352
rect 41140 74288 41204 74352
rect 41220 74288 41284 74352
rect 46740 74288 46804 74352
rect 46820 74288 46884 74352
rect 46900 74288 46964 74352
rect 46980 74288 47044 74352
rect 47060 74288 47124 74352
rect 47140 74288 47204 74352
rect 47220 74288 47284 74352
rect 52740 74288 52804 74352
rect 52820 74288 52884 74352
rect 52900 74288 52964 74352
rect 52980 74288 53044 74352
rect 53060 74288 53124 74352
rect 53140 74288 53204 74352
rect 53220 74288 53284 74352
rect 58740 74288 58804 74352
rect 58820 74288 58884 74352
rect 58900 74288 58964 74352
rect 58980 74288 59044 74352
rect 59060 74288 59124 74352
rect 59140 74288 59204 74352
rect 59220 74288 59284 74352
rect 64740 74288 64804 74352
rect 64820 74288 64884 74352
rect 64900 74288 64964 74352
rect 64980 74288 65044 74352
rect 65060 74288 65124 74352
rect 65140 74288 65204 74352
rect 65220 74288 65284 74352
rect 70740 74288 70804 74352
rect 70820 74288 70884 74352
rect 70900 74288 70964 74352
rect 70980 74288 71044 74352
rect 71060 74288 71124 74352
rect 71140 74288 71204 74352
rect 71220 74288 71284 74352
rect 1740 72176 1804 72240
rect 1820 72176 1884 72240
rect 1900 72176 1964 72240
rect 1980 72176 2044 72240
rect 2060 72176 2124 72240
rect 2140 72176 2204 72240
rect 2220 72176 2284 72240
rect 7740 72176 7804 72240
rect 7820 72176 7884 72240
rect 7900 72176 7964 72240
rect 7980 72176 8044 72240
rect 8060 72176 8124 72240
rect 8140 72176 8204 72240
rect 8220 72176 8284 72240
rect 13740 72176 13804 72240
rect 13820 72176 13884 72240
rect 13900 72176 13964 72240
rect 13980 72176 14044 72240
rect 14060 72176 14124 72240
rect 14140 72176 14204 72240
rect 14220 72176 14284 72240
rect 19740 72176 19804 72240
rect 19820 72176 19884 72240
rect 19900 72176 19964 72240
rect 19980 72176 20044 72240
rect 20060 72176 20124 72240
rect 20140 72176 20204 72240
rect 20220 72176 20284 72240
rect 25740 72176 25804 72240
rect 25820 72176 25884 72240
rect 25900 72176 25964 72240
rect 25980 72176 26044 72240
rect 26060 72176 26124 72240
rect 26140 72176 26204 72240
rect 26220 72176 26284 72240
rect 31740 72176 31804 72240
rect 31820 72176 31884 72240
rect 31900 72176 31964 72240
rect 31980 72176 32044 72240
rect 32060 72176 32124 72240
rect 32140 72176 32204 72240
rect 32220 72176 32284 72240
rect 37740 72176 37804 72240
rect 37820 72176 37884 72240
rect 37900 72176 37964 72240
rect 37980 72176 38044 72240
rect 38060 72176 38124 72240
rect 38140 72176 38204 72240
rect 38220 72176 38284 72240
rect 43740 72176 43804 72240
rect 43820 72176 43884 72240
rect 43900 72176 43964 72240
rect 43980 72176 44044 72240
rect 44060 72176 44124 72240
rect 44140 72176 44204 72240
rect 44220 72176 44284 72240
rect 49740 72176 49804 72240
rect 49820 72176 49884 72240
rect 49900 72176 49964 72240
rect 49980 72176 50044 72240
rect 50060 72176 50124 72240
rect 50140 72176 50204 72240
rect 50220 72176 50284 72240
rect 55740 72176 55804 72240
rect 55820 72176 55884 72240
rect 55900 72176 55964 72240
rect 55980 72176 56044 72240
rect 56060 72176 56124 72240
rect 56140 72176 56204 72240
rect 56220 72176 56284 72240
rect 61740 72176 61804 72240
rect 61820 72176 61884 72240
rect 61900 72176 61964 72240
rect 61980 72176 62044 72240
rect 62060 72176 62124 72240
rect 62140 72176 62204 72240
rect 62220 72176 62284 72240
rect 67740 72176 67804 72240
rect 67820 72176 67884 72240
rect 67900 72176 67964 72240
rect 67980 72176 68044 72240
rect 68060 72176 68124 72240
rect 68140 72176 68204 72240
rect 68220 72176 68284 72240
rect 73740 72176 73804 72240
rect 73820 72176 73884 72240
rect 73900 72176 73964 72240
rect 73980 72176 74044 72240
rect 74060 72176 74124 72240
rect 74140 72176 74204 72240
rect 74220 72176 74284 72240
rect 1740 72096 1804 72160
rect 1820 72096 1884 72160
rect 1900 72096 1964 72160
rect 1980 72096 2044 72160
rect 2060 72096 2124 72160
rect 2140 72096 2204 72160
rect 2220 72096 2284 72160
rect 7740 72096 7804 72160
rect 7820 72096 7884 72160
rect 7900 72096 7964 72160
rect 7980 72096 8044 72160
rect 8060 72096 8124 72160
rect 8140 72096 8204 72160
rect 8220 72096 8284 72160
rect 13740 72096 13804 72160
rect 13820 72096 13884 72160
rect 13900 72096 13964 72160
rect 13980 72096 14044 72160
rect 14060 72096 14124 72160
rect 14140 72096 14204 72160
rect 14220 72096 14284 72160
rect 19740 72096 19804 72160
rect 19820 72096 19884 72160
rect 19900 72096 19964 72160
rect 19980 72096 20044 72160
rect 20060 72096 20124 72160
rect 20140 72096 20204 72160
rect 20220 72096 20284 72160
rect 25740 72096 25804 72160
rect 25820 72096 25884 72160
rect 25900 72096 25964 72160
rect 25980 72096 26044 72160
rect 26060 72096 26124 72160
rect 26140 72096 26204 72160
rect 26220 72096 26284 72160
rect 31740 72096 31804 72160
rect 31820 72096 31884 72160
rect 31900 72096 31964 72160
rect 31980 72096 32044 72160
rect 32060 72096 32124 72160
rect 32140 72096 32204 72160
rect 32220 72096 32284 72160
rect 37740 72096 37804 72160
rect 37820 72096 37884 72160
rect 37900 72096 37964 72160
rect 37980 72096 38044 72160
rect 38060 72096 38124 72160
rect 38140 72096 38204 72160
rect 38220 72096 38284 72160
rect 43740 72096 43804 72160
rect 43820 72096 43884 72160
rect 43900 72096 43964 72160
rect 43980 72096 44044 72160
rect 44060 72096 44124 72160
rect 44140 72096 44204 72160
rect 44220 72096 44284 72160
rect 49740 72096 49804 72160
rect 49820 72096 49884 72160
rect 49900 72096 49964 72160
rect 49980 72096 50044 72160
rect 50060 72096 50124 72160
rect 50140 72096 50204 72160
rect 50220 72096 50284 72160
rect 55740 72096 55804 72160
rect 55820 72096 55884 72160
rect 55900 72096 55964 72160
rect 55980 72096 56044 72160
rect 56060 72096 56124 72160
rect 56140 72096 56204 72160
rect 56220 72096 56284 72160
rect 61740 72096 61804 72160
rect 61820 72096 61884 72160
rect 61900 72096 61964 72160
rect 61980 72096 62044 72160
rect 62060 72096 62124 72160
rect 62140 72096 62204 72160
rect 62220 72096 62284 72160
rect 67740 72096 67804 72160
rect 67820 72096 67884 72160
rect 67900 72096 67964 72160
rect 67980 72096 68044 72160
rect 68060 72096 68124 72160
rect 68140 72096 68204 72160
rect 68220 72096 68284 72160
rect 73740 72096 73804 72160
rect 73820 72096 73884 72160
rect 73900 72096 73964 72160
rect 73980 72096 74044 72160
rect 74060 72096 74124 72160
rect 74140 72096 74204 72160
rect 74220 72096 74284 72160
rect 1740 72016 1804 72080
rect 1820 72016 1884 72080
rect 1900 72016 1964 72080
rect 1980 72016 2044 72080
rect 2060 72016 2124 72080
rect 2140 72016 2204 72080
rect 2220 72016 2284 72080
rect 7740 72016 7804 72080
rect 7820 72016 7884 72080
rect 7900 72016 7964 72080
rect 7980 72016 8044 72080
rect 8060 72016 8124 72080
rect 8140 72016 8204 72080
rect 8220 72016 8284 72080
rect 13740 72016 13804 72080
rect 13820 72016 13884 72080
rect 13900 72016 13964 72080
rect 13980 72016 14044 72080
rect 14060 72016 14124 72080
rect 14140 72016 14204 72080
rect 14220 72016 14284 72080
rect 19740 72016 19804 72080
rect 19820 72016 19884 72080
rect 19900 72016 19964 72080
rect 19980 72016 20044 72080
rect 20060 72016 20124 72080
rect 20140 72016 20204 72080
rect 20220 72016 20284 72080
rect 25740 72016 25804 72080
rect 25820 72016 25884 72080
rect 25900 72016 25964 72080
rect 25980 72016 26044 72080
rect 26060 72016 26124 72080
rect 26140 72016 26204 72080
rect 26220 72016 26284 72080
rect 31740 72016 31804 72080
rect 31820 72016 31884 72080
rect 31900 72016 31964 72080
rect 31980 72016 32044 72080
rect 32060 72016 32124 72080
rect 32140 72016 32204 72080
rect 32220 72016 32284 72080
rect 37740 72016 37804 72080
rect 37820 72016 37884 72080
rect 37900 72016 37964 72080
rect 37980 72016 38044 72080
rect 38060 72016 38124 72080
rect 38140 72016 38204 72080
rect 38220 72016 38284 72080
rect 43740 72016 43804 72080
rect 43820 72016 43884 72080
rect 43900 72016 43964 72080
rect 43980 72016 44044 72080
rect 44060 72016 44124 72080
rect 44140 72016 44204 72080
rect 44220 72016 44284 72080
rect 49740 72016 49804 72080
rect 49820 72016 49884 72080
rect 49900 72016 49964 72080
rect 49980 72016 50044 72080
rect 50060 72016 50124 72080
rect 50140 72016 50204 72080
rect 50220 72016 50284 72080
rect 55740 72016 55804 72080
rect 55820 72016 55884 72080
rect 55900 72016 55964 72080
rect 55980 72016 56044 72080
rect 56060 72016 56124 72080
rect 56140 72016 56204 72080
rect 56220 72016 56284 72080
rect 61740 72016 61804 72080
rect 61820 72016 61884 72080
rect 61900 72016 61964 72080
rect 61980 72016 62044 72080
rect 62060 72016 62124 72080
rect 62140 72016 62204 72080
rect 62220 72016 62284 72080
rect 67740 72016 67804 72080
rect 67820 72016 67884 72080
rect 67900 72016 67964 72080
rect 67980 72016 68044 72080
rect 68060 72016 68124 72080
rect 68140 72016 68204 72080
rect 68220 72016 68284 72080
rect 73740 72016 73804 72080
rect 73820 72016 73884 72080
rect 73900 72016 73964 72080
rect 73980 72016 74044 72080
rect 74060 72016 74124 72080
rect 74140 72016 74204 72080
rect 74220 72016 74284 72080
rect 1740 71936 1804 72000
rect 1820 71936 1884 72000
rect 1900 71936 1964 72000
rect 1980 71936 2044 72000
rect 2060 71936 2124 72000
rect 2140 71936 2204 72000
rect 2220 71936 2284 72000
rect 7740 71936 7804 72000
rect 7820 71936 7884 72000
rect 7900 71936 7964 72000
rect 7980 71936 8044 72000
rect 8060 71936 8124 72000
rect 8140 71936 8204 72000
rect 8220 71936 8284 72000
rect 13740 71936 13804 72000
rect 13820 71936 13884 72000
rect 13900 71936 13964 72000
rect 13980 71936 14044 72000
rect 14060 71936 14124 72000
rect 14140 71936 14204 72000
rect 14220 71936 14284 72000
rect 19740 71936 19804 72000
rect 19820 71936 19884 72000
rect 19900 71936 19964 72000
rect 19980 71936 20044 72000
rect 20060 71936 20124 72000
rect 20140 71936 20204 72000
rect 20220 71936 20284 72000
rect 25740 71936 25804 72000
rect 25820 71936 25884 72000
rect 25900 71936 25964 72000
rect 25980 71936 26044 72000
rect 26060 71936 26124 72000
rect 26140 71936 26204 72000
rect 26220 71936 26284 72000
rect 31740 71936 31804 72000
rect 31820 71936 31884 72000
rect 31900 71936 31964 72000
rect 31980 71936 32044 72000
rect 32060 71936 32124 72000
rect 32140 71936 32204 72000
rect 32220 71936 32284 72000
rect 37740 71936 37804 72000
rect 37820 71936 37884 72000
rect 37900 71936 37964 72000
rect 37980 71936 38044 72000
rect 38060 71936 38124 72000
rect 38140 71936 38204 72000
rect 38220 71936 38284 72000
rect 43740 71936 43804 72000
rect 43820 71936 43884 72000
rect 43900 71936 43964 72000
rect 43980 71936 44044 72000
rect 44060 71936 44124 72000
rect 44140 71936 44204 72000
rect 44220 71936 44284 72000
rect 49740 71936 49804 72000
rect 49820 71936 49884 72000
rect 49900 71936 49964 72000
rect 49980 71936 50044 72000
rect 50060 71936 50124 72000
rect 50140 71936 50204 72000
rect 50220 71936 50284 72000
rect 55740 71936 55804 72000
rect 55820 71936 55884 72000
rect 55900 71936 55964 72000
rect 55980 71936 56044 72000
rect 56060 71936 56124 72000
rect 56140 71936 56204 72000
rect 56220 71936 56284 72000
rect 61740 71936 61804 72000
rect 61820 71936 61884 72000
rect 61900 71936 61964 72000
rect 61980 71936 62044 72000
rect 62060 71936 62124 72000
rect 62140 71936 62204 72000
rect 62220 71936 62284 72000
rect 67740 71936 67804 72000
rect 67820 71936 67884 72000
rect 67900 71936 67964 72000
rect 67980 71936 68044 72000
rect 68060 71936 68124 72000
rect 68140 71936 68204 72000
rect 68220 71936 68284 72000
rect 73740 71936 73804 72000
rect 73820 71936 73884 72000
rect 73900 71936 73964 72000
rect 73980 71936 74044 72000
rect 74060 71936 74124 72000
rect 74140 71936 74204 72000
rect 74220 71936 74284 72000
rect 4740 64528 4804 64592
rect 4820 64528 4884 64592
rect 4900 64528 4964 64592
rect 4980 64528 5044 64592
rect 5060 64528 5124 64592
rect 5140 64528 5204 64592
rect 5220 64528 5284 64592
rect 10740 64528 10804 64592
rect 10820 64528 10884 64592
rect 10900 64528 10964 64592
rect 10980 64528 11044 64592
rect 11060 64528 11124 64592
rect 11140 64528 11204 64592
rect 11220 64528 11284 64592
rect 16740 64528 16804 64592
rect 16820 64528 16884 64592
rect 16900 64528 16964 64592
rect 16980 64528 17044 64592
rect 17060 64528 17124 64592
rect 17140 64528 17204 64592
rect 17220 64528 17284 64592
rect 22740 64528 22804 64592
rect 22820 64528 22884 64592
rect 22900 64528 22964 64592
rect 22980 64528 23044 64592
rect 23060 64528 23124 64592
rect 23140 64528 23204 64592
rect 23220 64528 23284 64592
rect 28740 64528 28804 64592
rect 28820 64528 28884 64592
rect 28900 64528 28964 64592
rect 28980 64528 29044 64592
rect 29060 64528 29124 64592
rect 29140 64528 29204 64592
rect 29220 64528 29284 64592
rect 34740 64528 34804 64592
rect 34820 64528 34884 64592
rect 34900 64528 34964 64592
rect 34980 64528 35044 64592
rect 35060 64528 35124 64592
rect 35140 64528 35204 64592
rect 35220 64528 35284 64592
rect 40740 64528 40804 64592
rect 40820 64528 40884 64592
rect 40900 64528 40964 64592
rect 40980 64528 41044 64592
rect 41060 64528 41124 64592
rect 41140 64528 41204 64592
rect 41220 64528 41284 64592
rect 46740 64528 46804 64592
rect 46820 64528 46884 64592
rect 46900 64528 46964 64592
rect 46980 64528 47044 64592
rect 47060 64528 47124 64592
rect 47140 64528 47204 64592
rect 47220 64528 47284 64592
rect 52740 64528 52804 64592
rect 52820 64528 52884 64592
rect 52900 64528 52964 64592
rect 52980 64528 53044 64592
rect 53060 64528 53124 64592
rect 53140 64528 53204 64592
rect 53220 64528 53284 64592
rect 58740 64528 58804 64592
rect 58820 64528 58884 64592
rect 58900 64528 58964 64592
rect 58980 64528 59044 64592
rect 59060 64528 59124 64592
rect 59140 64528 59204 64592
rect 59220 64528 59284 64592
rect 64740 64528 64804 64592
rect 64820 64528 64884 64592
rect 64900 64528 64964 64592
rect 64980 64528 65044 64592
rect 65060 64528 65124 64592
rect 65140 64528 65204 64592
rect 65220 64528 65284 64592
rect 70740 64528 70804 64592
rect 70820 64528 70884 64592
rect 70900 64528 70964 64592
rect 70980 64528 71044 64592
rect 71060 64528 71124 64592
rect 71140 64528 71204 64592
rect 71220 64528 71284 64592
rect 4740 64448 4804 64512
rect 4820 64448 4884 64512
rect 4900 64448 4964 64512
rect 4980 64448 5044 64512
rect 5060 64448 5124 64512
rect 5140 64448 5204 64512
rect 5220 64448 5284 64512
rect 10740 64448 10804 64512
rect 10820 64448 10884 64512
rect 10900 64448 10964 64512
rect 10980 64448 11044 64512
rect 11060 64448 11124 64512
rect 11140 64448 11204 64512
rect 11220 64448 11284 64512
rect 16740 64448 16804 64512
rect 16820 64448 16884 64512
rect 16900 64448 16964 64512
rect 16980 64448 17044 64512
rect 17060 64448 17124 64512
rect 17140 64448 17204 64512
rect 17220 64448 17284 64512
rect 22740 64448 22804 64512
rect 22820 64448 22884 64512
rect 22900 64448 22964 64512
rect 22980 64448 23044 64512
rect 23060 64448 23124 64512
rect 23140 64448 23204 64512
rect 23220 64448 23284 64512
rect 28740 64448 28804 64512
rect 28820 64448 28884 64512
rect 28900 64448 28964 64512
rect 28980 64448 29044 64512
rect 29060 64448 29124 64512
rect 29140 64448 29204 64512
rect 29220 64448 29284 64512
rect 34740 64448 34804 64512
rect 34820 64448 34884 64512
rect 34900 64448 34964 64512
rect 34980 64448 35044 64512
rect 35060 64448 35124 64512
rect 35140 64448 35204 64512
rect 35220 64448 35284 64512
rect 40740 64448 40804 64512
rect 40820 64448 40884 64512
rect 40900 64448 40964 64512
rect 40980 64448 41044 64512
rect 41060 64448 41124 64512
rect 41140 64448 41204 64512
rect 41220 64448 41284 64512
rect 46740 64448 46804 64512
rect 46820 64448 46884 64512
rect 46900 64448 46964 64512
rect 46980 64448 47044 64512
rect 47060 64448 47124 64512
rect 47140 64448 47204 64512
rect 47220 64448 47284 64512
rect 52740 64448 52804 64512
rect 52820 64448 52884 64512
rect 52900 64448 52964 64512
rect 52980 64448 53044 64512
rect 53060 64448 53124 64512
rect 53140 64448 53204 64512
rect 53220 64448 53284 64512
rect 58740 64448 58804 64512
rect 58820 64448 58884 64512
rect 58900 64448 58964 64512
rect 58980 64448 59044 64512
rect 59060 64448 59124 64512
rect 59140 64448 59204 64512
rect 59220 64448 59284 64512
rect 64740 64448 64804 64512
rect 64820 64448 64884 64512
rect 64900 64448 64964 64512
rect 64980 64448 65044 64512
rect 65060 64448 65124 64512
rect 65140 64448 65204 64512
rect 65220 64448 65284 64512
rect 70740 64448 70804 64512
rect 70820 64448 70884 64512
rect 70900 64448 70964 64512
rect 70980 64448 71044 64512
rect 71060 64448 71124 64512
rect 71140 64448 71204 64512
rect 71220 64448 71284 64512
rect 4740 64368 4804 64432
rect 4820 64368 4884 64432
rect 4900 64368 4964 64432
rect 4980 64368 5044 64432
rect 5060 64368 5124 64432
rect 5140 64368 5204 64432
rect 5220 64368 5284 64432
rect 10740 64368 10804 64432
rect 10820 64368 10884 64432
rect 10900 64368 10964 64432
rect 10980 64368 11044 64432
rect 11060 64368 11124 64432
rect 11140 64368 11204 64432
rect 11220 64368 11284 64432
rect 16740 64368 16804 64432
rect 16820 64368 16884 64432
rect 16900 64368 16964 64432
rect 16980 64368 17044 64432
rect 17060 64368 17124 64432
rect 17140 64368 17204 64432
rect 17220 64368 17284 64432
rect 22740 64368 22804 64432
rect 22820 64368 22884 64432
rect 22900 64368 22964 64432
rect 22980 64368 23044 64432
rect 23060 64368 23124 64432
rect 23140 64368 23204 64432
rect 23220 64368 23284 64432
rect 28740 64368 28804 64432
rect 28820 64368 28884 64432
rect 28900 64368 28964 64432
rect 28980 64368 29044 64432
rect 29060 64368 29124 64432
rect 29140 64368 29204 64432
rect 29220 64368 29284 64432
rect 34740 64368 34804 64432
rect 34820 64368 34884 64432
rect 34900 64368 34964 64432
rect 34980 64368 35044 64432
rect 35060 64368 35124 64432
rect 35140 64368 35204 64432
rect 35220 64368 35284 64432
rect 40740 64368 40804 64432
rect 40820 64368 40884 64432
rect 40900 64368 40964 64432
rect 40980 64368 41044 64432
rect 41060 64368 41124 64432
rect 41140 64368 41204 64432
rect 41220 64368 41284 64432
rect 46740 64368 46804 64432
rect 46820 64368 46884 64432
rect 46900 64368 46964 64432
rect 46980 64368 47044 64432
rect 47060 64368 47124 64432
rect 47140 64368 47204 64432
rect 47220 64368 47284 64432
rect 52740 64368 52804 64432
rect 52820 64368 52884 64432
rect 52900 64368 52964 64432
rect 52980 64368 53044 64432
rect 53060 64368 53124 64432
rect 53140 64368 53204 64432
rect 53220 64368 53284 64432
rect 58740 64368 58804 64432
rect 58820 64368 58884 64432
rect 58900 64368 58964 64432
rect 58980 64368 59044 64432
rect 59060 64368 59124 64432
rect 59140 64368 59204 64432
rect 59220 64368 59284 64432
rect 64740 64368 64804 64432
rect 64820 64368 64884 64432
rect 64900 64368 64964 64432
rect 64980 64368 65044 64432
rect 65060 64368 65124 64432
rect 65140 64368 65204 64432
rect 65220 64368 65284 64432
rect 70740 64368 70804 64432
rect 70820 64368 70884 64432
rect 70900 64368 70964 64432
rect 70980 64368 71044 64432
rect 71060 64368 71124 64432
rect 71140 64368 71204 64432
rect 71220 64368 71284 64432
rect 4740 64288 4804 64352
rect 4820 64288 4884 64352
rect 4900 64288 4964 64352
rect 4980 64288 5044 64352
rect 5060 64288 5124 64352
rect 5140 64288 5204 64352
rect 5220 64288 5284 64352
rect 10740 64288 10804 64352
rect 10820 64288 10884 64352
rect 10900 64288 10964 64352
rect 10980 64288 11044 64352
rect 11060 64288 11124 64352
rect 11140 64288 11204 64352
rect 11220 64288 11284 64352
rect 16740 64288 16804 64352
rect 16820 64288 16884 64352
rect 16900 64288 16964 64352
rect 16980 64288 17044 64352
rect 17060 64288 17124 64352
rect 17140 64288 17204 64352
rect 17220 64288 17284 64352
rect 22740 64288 22804 64352
rect 22820 64288 22884 64352
rect 22900 64288 22964 64352
rect 22980 64288 23044 64352
rect 23060 64288 23124 64352
rect 23140 64288 23204 64352
rect 23220 64288 23284 64352
rect 28740 64288 28804 64352
rect 28820 64288 28884 64352
rect 28900 64288 28964 64352
rect 28980 64288 29044 64352
rect 29060 64288 29124 64352
rect 29140 64288 29204 64352
rect 29220 64288 29284 64352
rect 34740 64288 34804 64352
rect 34820 64288 34884 64352
rect 34900 64288 34964 64352
rect 34980 64288 35044 64352
rect 35060 64288 35124 64352
rect 35140 64288 35204 64352
rect 35220 64288 35284 64352
rect 40740 64288 40804 64352
rect 40820 64288 40884 64352
rect 40900 64288 40964 64352
rect 40980 64288 41044 64352
rect 41060 64288 41124 64352
rect 41140 64288 41204 64352
rect 41220 64288 41284 64352
rect 46740 64288 46804 64352
rect 46820 64288 46884 64352
rect 46900 64288 46964 64352
rect 46980 64288 47044 64352
rect 47060 64288 47124 64352
rect 47140 64288 47204 64352
rect 47220 64288 47284 64352
rect 52740 64288 52804 64352
rect 52820 64288 52884 64352
rect 52900 64288 52964 64352
rect 52980 64288 53044 64352
rect 53060 64288 53124 64352
rect 53140 64288 53204 64352
rect 53220 64288 53284 64352
rect 58740 64288 58804 64352
rect 58820 64288 58884 64352
rect 58900 64288 58964 64352
rect 58980 64288 59044 64352
rect 59060 64288 59124 64352
rect 59140 64288 59204 64352
rect 59220 64288 59284 64352
rect 64740 64288 64804 64352
rect 64820 64288 64884 64352
rect 64900 64288 64964 64352
rect 64980 64288 65044 64352
rect 65060 64288 65124 64352
rect 65140 64288 65204 64352
rect 65220 64288 65284 64352
rect 70740 64288 70804 64352
rect 70820 64288 70884 64352
rect 70900 64288 70964 64352
rect 70980 64288 71044 64352
rect 71060 64288 71124 64352
rect 71140 64288 71204 64352
rect 71220 64288 71284 64352
rect 1740 62176 1804 62240
rect 1820 62176 1884 62240
rect 1900 62176 1964 62240
rect 1980 62176 2044 62240
rect 2060 62176 2124 62240
rect 2140 62176 2204 62240
rect 2220 62176 2284 62240
rect 7740 62176 7804 62240
rect 7820 62176 7884 62240
rect 7900 62176 7964 62240
rect 7980 62176 8044 62240
rect 8060 62176 8124 62240
rect 8140 62176 8204 62240
rect 8220 62176 8284 62240
rect 13740 62176 13804 62240
rect 13820 62176 13884 62240
rect 13900 62176 13964 62240
rect 13980 62176 14044 62240
rect 14060 62176 14124 62240
rect 14140 62176 14204 62240
rect 14220 62176 14284 62240
rect 19740 62176 19804 62240
rect 19820 62176 19884 62240
rect 19900 62176 19964 62240
rect 19980 62176 20044 62240
rect 20060 62176 20124 62240
rect 20140 62176 20204 62240
rect 20220 62176 20284 62240
rect 25740 62176 25804 62240
rect 25820 62176 25884 62240
rect 25900 62176 25964 62240
rect 25980 62176 26044 62240
rect 26060 62176 26124 62240
rect 26140 62176 26204 62240
rect 26220 62176 26284 62240
rect 31740 62176 31804 62240
rect 31820 62176 31884 62240
rect 31900 62176 31964 62240
rect 31980 62176 32044 62240
rect 32060 62176 32124 62240
rect 32140 62176 32204 62240
rect 32220 62176 32284 62240
rect 37740 62176 37804 62240
rect 37820 62176 37884 62240
rect 37900 62176 37964 62240
rect 37980 62176 38044 62240
rect 38060 62176 38124 62240
rect 38140 62176 38204 62240
rect 38220 62176 38284 62240
rect 43740 62176 43804 62240
rect 43820 62176 43884 62240
rect 43900 62176 43964 62240
rect 43980 62176 44044 62240
rect 44060 62176 44124 62240
rect 44140 62176 44204 62240
rect 44220 62176 44284 62240
rect 49740 62176 49804 62240
rect 49820 62176 49884 62240
rect 49900 62176 49964 62240
rect 49980 62176 50044 62240
rect 50060 62176 50124 62240
rect 50140 62176 50204 62240
rect 50220 62176 50284 62240
rect 55740 62176 55804 62240
rect 55820 62176 55884 62240
rect 55900 62176 55964 62240
rect 55980 62176 56044 62240
rect 56060 62176 56124 62240
rect 56140 62176 56204 62240
rect 56220 62176 56284 62240
rect 61740 62176 61804 62240
rect 61820 62176 61884 62240
rect 61900 62176 61964 62240
rect 61980 62176 62044 62240
rect 62060 62176 62124 62240
rect 62140 62176 62204 62240
rect 62220 62176 62284 62240
rect 67740 62176 67804 62240
rect 67820 62176 67884 62240
rect 67900 62176 67964 62240
rect 67980 62176 68044 62240
rect 68060 62176 68124 62240
rect 68140 62176 68204 62240
rect 68220 62176 68284 62240
rect 73740 62176 73804 62240
rect 73820 62176 73884 62240
rect 73900 62176 73964 62240
rect 73980 62176 74044 62240
rect 74060 62176 74124 62240
rect 74140 62176 74204 62240
rect 74220 62176 74284 62240
rect 1740 62096 1804 62160
rect 1820 62096 1884 62160
rect 1900 62096 1964 62160
rect 1980 62096 2044 62160
rect 2060 62096 2124 62160
rect 2140 62096 2204 62160
rect 2220 62096 2284 62160
rect 7740 62096 7804 62160
rect 7820 62096 7884 62160
rect 7900 62096 7964 62160
rect 7980 62096 8044 62160
rect 8060 62096 8124 62160
rect 8140 62096 8204 62160
rect 8220 62096 8284 62160
rect 13740 62096 13804 62160
rect 13820 62096 13884 62160
rect 13900 62096 13964 62160
rect 13980 62096 14044 62160
rect 14060 62096 14124 62160
rect 14140 62096 14204 62160
rect 14220 62096 14284 62160
rect 19740 62096 19804 62160
rect 19820 62096 19884 62160
rect 19900 62096 19964 62160
rect 19980 62096 20044 62160
rect 20060 62096 20124 62160
rect 20140 62096 20204 62160
rect 20220 62096 20284 62160
rect 25740 62096 25804 62160
rect 25820 62096 25884 62160
rect 25900 62096 25964 62160
rect 25980 62096 26044 62160
rect 26060 62096 26124 62160
rect 26140 62096 26204 62160
rect 26220 62096 26284 62160
rect 31740 62096 31804 62160
rect 31820 62096 31884 62160
rect 31900 62096 31964 62160
rect 31980 62096 32044 62160
rect 32060 62096 32124 62160
rect 32140 62096 32204 62160
rect 32220 62096 32284 62160
rect 37740 62096 37804 62160
rect 37820 62096 37884 62160
rect 37900 62096 37964 62160
rect 37980 62096 38044 62160
rect 38060 62096 38124 62160
rect 38140 62096 38204 62160
rect 38220 62096 38284 62160
rect 43740 62096 43804 62160
rect 43820 62096 43884 62160
rect 43900 62096 43964 62160
rect 43980 62096 44044 62160
rect 44060 62096 44124 62160
rect 44140 62096 44204 62160
rect 44220 62096 44284 62160
rect 49740 62096 49804 62160
rect 49820 62096 49884 62160
rect 49900 62096 49964 62160
rect 49980 62096 50044 62160
rect 50060 62096 50124 62160
rect 50140 62096 50204 62160
rect 50220 62096 50284 62160
rect 55740 62096 55804 62160
rect 55820 62096 55884 62160
rect 55900 62096 55964 62160
rect 55980 62096 56044 62160
rect 56060 62096 56124 62160
rect 56140 62096 56204 62160
rect 56220 62096 56284 62160
rect 61740 62096 61804 62160
rect 61820 62096 61884 62160
rect 61900 62096 61964 62160
rect 61980 62096 62044 62160
rect 62060 62096 62124 62160
rect 62140 62096 62204 62160
rect 62220 62096 62284 62160
rect 67740 62096 67804 62160
rect 67820 62096 67884 62160
rect 67900 62096 67964 62160
rect 67980 62096 68044 62160
rect 68060 62096 68124 62160
rect 68140 62096 68204 62160
rect 68220 62096 68284 62160
rect 73740 62096 73804 62160
rect 73820 62096 73884 62160
rect 73900 62096 73964 62160
rect 73980 62096 74044 62160
rect 74060 62096 74124 62160
rect 74140 62096 74204 62160
rect 74220 62096 74284 62160
rect 1740 62016 1804 62080
rect 1820 62016 1884 62080
rect 1900 62016 1964 62080
rect 1980 62016 2044 62080
rect 2060 62016 2124 62080
rect 2140 62016 2204 62080
rect 2220 62016 2284 62080
rect 7740 62016 7804 62080
rect 7820 62016 7884 62080
rect 7900 62016 7964 62080
rect 7980 62016 8044 62080
rect 8060 62016 8124 62080
rect 8140 62016 8204 62080
rect 8220 62016 8284 62080
rect 13740 62016 13804 62080
rect 13820 62016 13884 62080
rect 13900 62016 13964 62080
rect 13980 62016 14044 62080
rect 14060 62016 14124 62080
rect 14140 62016 14204 62080
rect 14220 62016 14284 62080
rect 19740 62016 19804 62080
rect 19820 62016 19884 62080
rect 19900 62016 19964 62080
rect 19980 62016 20044 62080
rect 20060 62016 20124 62080
rect 20140 62016 20204 62080
rect 20220 62016 20284 62080
rect 25740 62016 25804 62080
rect 25820 62016 25884 62080
rect 25900 62016 25964 62080
rect 25980 62016 26044 62080
rect 26060 62016 26124 62080
rect 26140 62016 26204 62080
rect 26220 62016 26284 62080
rect 31740 62016 31804 62080
rect 31820 62016 31884 62080
rect 31900 62016 31964 62080
rect 31980 62016 32044 62080
rect 32060 62016 32124 62080
rect 32140 62016 32204 62080
rect 32220 62016 32284 62080
rect 37740 62016 37804 62080
rect 37820 62016 37884 62080
rect 37900 62016 37964 62080
rect 37980 62016 38044 62080
rect 38060 62016 38124 62080
rect 38140 62016 38204 62080
rect 38220 62016 38284 62080
rect 43740 62016 43804 62080
rect 43820 62016 43884 62080
rect 43900 62016 43964 62080
rect 43980 62016 44044 62080
rect 44060 62016 44124 62080
rect 44140 62016 44204 62080
rect 44220 62016 44284 62080
rect 49740 62016 49804 62080
rect 49820 62016 49884 62080
rect 49900 62016 49964 62080
rect 49980 62016 50044 62080
rect 50060 62016 50124 62080
rect 50140 62016 50204 62080
rect 50220 62016 50284 62080
rect 55740 62016 55804 62080
rect 55820 62016 55884 62080
rect 55900 62016 55964 62080
rect 55980 62016 56044 62080
rect 56060 62016 56124 62080
rect 56140 62016 56204 62080
rect 56220 62016 56284 62080
rect 61740 62016 61804 62080
rect 61820 62016 61884 62080
rect 61900 62016 61964 62080
rect 61980 62016 62044 62080
rect 62060 62016 62124 62080
rect 62140 62016 62204 62080
rect 62220 62016 62284 62080
rect 67740 62016 67804 62080
rect 67820 62016 67884 62080
rect 67900 62016 67964 62080
rect 67980 62016 68044 62080
rect 68060 62016 68124 62080
rect 68140 62016 68204 62080
rect 68220 62016 68284 62080
rect 73740 62016 73804 62080
rect 73820 62016 73884 62080
rect 73900 62016 73964 62080
rect 73980 62016 74044 62080
rect 74060 62016 74124 62080
rect 74140 62016 74204 62080
rect 74220 62016 74284 62080
rect 1740 61936 1804 62000
rect 1820 61936 1884 62000
rect 1900 61936 1964 62000
rect 1980 61936 2044 62000
rect 2060 61936 2124 62000
rect 2140 61936 2204 62000
rect 2220 61936 2284 62000
rect 7740 61936 7804 62000
rect 7820 61936 7884 62000
rect 7900 61936 7964 62000
rect 7980 61936 8044 62000
rect 8060 61936 8124 62000
rect 8140 61936 8204 62000
rect 8220 61936 8284 62000
rect 13740 61936 13804 62000
rect 13820 61936 13884 62000
rect 13900 61936 13964 62000
rect 13980 61936 14044 62000
rect 14060 61936 14124 62000
rect 14140 61936 14204 62000
rect 14220 61936 14284 62000
rect 19740 61936 19804 62000
rect 19820 61936 19884 62000
rect 19900 61936 19964 62000
rect 19980 61936 20044 62000
rect 20060 61936 20124 62000
rect 20140 61936 20204 62000
rect 20220 61936 20284 62000
rect 25740 61936 25804 62000
rect 25820 61936 25884 62000
rect 25900 61936 25964 62000
rect 25980 61936 26044 62000
rect 26060 61936 26124 62000
rect 26140 61936 26204 62000
rect 26220 61936 26284 62000
rect 31740 61936 31804 62000
rect 31820 61936 31884 62000
rect 31900 61936 31964 62000
rect 31980 61936 32044 62000
rect 32060 61936 32124 62000
rect 32140 61936 32204 62000
rect 32220 61936 32284 62000
rect 37740 61936 37804 62000
rect 37820 61936 37884 62000
rect 37900 61936 37964 62000
rect 37980 61936 38044 62000
rect 38060 61936 38124 62000
rect 38140 61936 38204 62000
rect 38220 61936 38284 62000
rect 43740 61936 43804 62000
rect 43820 61936 43884 62000
rect 43900 61936 43964 62000
rect 43980 61936 44044 62000
rect 44060 61936 44124 62000
rect 44140 61936 44204 62000
rect 44220 61936 44284 62000
rect 49740 61936 49804 62000
rect 49820 61936 49884 62000
rect 49900 61936 49964 62000
rect 49980 61936 50044 62000
rect 50060 61936 50124 62000
rect 50140 61936 50204 62000
rect 50220 61936 50284 62000
rect 55740 61936 55804 62000
rect 55820 61936 55884 62000
rect 55900 61936 55964 62000
rect 55980 61936 56044 62000
rect 56060 61936 56124 62000
rect 56140 61936 56204 62000
rect 56220 61936 56284 62000
rect 61740 61936 61804 62000
rect 61820 61936 61884 62000
rect 61900 61936 61964 62000
rect 61980 61936 62044 62000
rect 62060 61936 62124 62000
rect 62140 61936 62204 62000
rect 62220 61936 62284 62000
rect 67740 61936 67804 62000
rect 67820 61936 67884 62000
rect 67900 61936 67964 62000
rect 67980 61936 68044 62000
rect 68060 61936 68124 62000
rect 68140 61936 68204 62000
rect 68220 61936 68284 62000
rect 73740 61936 73804 62000
rect 73820 61936 73884 62000
rect 73900 61936 73964 62000
rect 73980 61936 74044 62000
rect 74060 61936 74124 62000
rect 74140 61936 74204 62000
rect 74220 61936 74284 62000
rect 4740 54528 4804 54592
rect 4820 54528 4884 54592
rect 4900 54528 4964 54592
rect 4980 54528 5044 54592
rect 5060 54528 5124 54592
rect 5140 54528 5204 54592
rect 5220 54528 5284 54592
rect 10740 54528 10804 54592
rect 10820 54528 10884 54592
rect 10900 54528 10964 54592
rect 10980 54528 11044 54592
rect 11060 54528 11124 54592
rect 11140 54528 11204 54592
rect 11220 54528 11284 54592
rect 16740 54528 16804 54592
rect 16820 54528 16884 54592
rect 16900 54528 16964 54592
rect 16980 54528 17044 54592
rect 17060 54528 17124 54592
rect 17140 54528 17204 54592
rect 17220 54528 17284 54592
rect 22740 54528 22804 54592
rect 22820 54528 22884 54592
rect 22900 54528 22964 54592
rect 22980 54528 23044 54592
rect 23060 54528 23124 54592
rect 23140 54528 23204 54592
rect 23220 54528 23284 54592
rect 28740 54528 28804 54592
rect 28820 54528 28884 54592
rect 28900 54528 28964 54592
rect 28980 54528 29044 54592
rect 29060 54528 29124 54592
rect 29140 54528 29204 54592
rect 29220 54528 29284 54592
rect 34740 54528 34804 54592
rect 34820 54528 34884 54592
rect 34900 54528 34964 54592
rect 34980 54528 35044 54592
rect 35060 54528 35124 54592
rect 35140 54528 35204 54592
rect 35220 54528 35284 54592
rect 40740 54528 40804 54592
rect 40820 54528 40884 54592
rect 40900 54528 40964 54592
rect 40980 54528 41044 54592
rect 41060 54528 41124 54592
rect 41140 54528 41204 54592
rect 41220 54528 41284 54592
rect 46740 54528 46804 54592
rect 46820 54528 46884 54592
rect 46900 54528 46964 54592
rect 46980 54528 47044 54592
rect 47060 54528 47124 54592
rect 47140 54528 47204 54592
rect 47220 54528 47284 54592
rect 52740 54528 52804 54592
rect 52820 54528 52884 54592
rect 52900 54528 52964 54592
rect 52980 54528 53044 54592
rect 53060 54528 53124 54592
rect 53140 54528 53204 54592
rect 53220 54528 53284 54592
rect 58740 54528 58804 54592
rect 58820 54528 58884 54592
rect 58900 54528 58964 54592
rect 58980 54528 59044 54592
rect 59060 54528 59124 54592
rect 59140 54528 59204 54592
rect 59220 54528 59284 54592
rect 64740 54528 64804 54592
rect 64820 54528 64884 54592
rect 64900 54528 64964 54592
rect 64980 54528 65044 54592
rect 65060 54528 65124 54592
rect 65140 54528 65204 54592
rect 65220 54528 65284 54592
rect 70740 54528 70804 54592
rect 70820 54528 70884 54592
rect 70900 54528 70964 54592
rect 70980 54528 71044 54592
rect 71060 54528 71124 54592
rect 71140 54528 71204 54592
rect 71220 54528 71284 54592
rect 4740 54448 4804 54512
rect 4820 54448 4884 54512
rect 4900 54448 4964 54512
rect 4980 54448 5044 54512
rect 5060 54448 5124 54512
rect 5140 54448 5204 54512
rect 5220 54448 5284 54512
rect 10740 54448 10804 54512
rect 10820 54448 10884 54512
rect 10900 54448 10964 54512
rect 10980 54448 11044 54512
rect 11060 54448 11124 54512
rect 11140 54448 11204 54512
rect 11220 54448 11284 54512
rect 16740 54448 16804 54512
rect 16820 54448 16884 54512
rect 16900 54448 16964 54512
rect 16980 54448 17044 54512
rect 17060 54448 17124 54512
rect 17140 54448 17204 54512
rect 17220 54448 17284 54512
rect 22740 54448 22804 54512
rect 22820 54448 22884 54512
rect 22900 54448 22964 54512
rect 22980 54448 23044 54512
rect 23060 54448 23124 54512
rect 23140 54448 23204 54512
rect 23220 54448 23284 54512
rect 28740 54448 28804 54512
rect 28820 54448 28884 54512
rect 28900 54448 28964 54512
rect 28980 54448 29044 54512
rect 29060 54448 29124 54512
rect 29140 54448 29204 54512
rect 29220 54448 29284 54512
rect 34740 54448 34804 54512
rect 34820 54448 34884 54512
rect 34900 54448 34964 54512
rect 34980 54448 35044 54512
rect 35060 54448 35124 54512
rect 35140 54448 35204 54512
rect 35220 54448 35284 54512
rect 40740 54448 40804 54512
rect 40820 54448 40884 54512
rect 40900 54448 40964 54512
rect 40980 54448 41044 54512
rect 41060 54448 41124 54512
rect 41140 54448 41204 54512
rect 41220 54448 41284 54512
rect 46740 54448 46804 54512
rect 46820 54448 46884 54512
rect 46900 54448 46964 54512
rect 46980 54448 47044 54512
rect 47060 54448 47124 54512
rect 47140 54448 47204 54512
rect 47220 54448 47284 54512
rect 52740 54448 52804 54512
rect 52820 54448 52884 54512
rect 52900 54448 52964 54512
rect 52980 54448 53044 54512
rect 53060 54448 53124 54512
rect 53140 54448 53204 54512
rect 53220 54448 53284 54512
rect 58740 54448 58804 54512
rect 58820 54448 58884 54512
rect 58900 54448 58964 54512
rect 58980 54448 59044 54512
rect 59060 54448 59124 54512
rect 59140 54448 59204 54512
rect 59220 54448 59284 54512
rect 64740 54448 64804 54512
rect 64820 54448 64884 54512
rect 64900 54448 64964 54512
rect 64980 54448 65044 54512
rect 65060 54448 65124 54512
rect 65140 54448 65204 54512
rect 65220 54448 65284 54512
rect 70740 54448 70804 54512
rect 70820 54448 70884 54512
rect 70900 54448 70964 54512
rect 70980 54448 71044 54512
rect 71060 54448 71124 54512
rect 71140 54448 71204 54512
rect 71220 54448 71284 54512
rect 4740 54368 4804 54432
rect 4820 54368 4884 54432
rect 4900 54368 4964 54432
rect 4980 54368 5044 54432
rect 5060 54368 5124 54432
rect 5140 54368 5204 54432
rect 5220 54368 5284 54432
rect 10740 54368 10804 54432
rect 10820 54368 10884 54432
rect 10900 54368 10964 54432
rect 10980 54368 11044 54432
rect 11060 54368 11124 54432
rect 11140 54368 11204 54432
rect 11220 54368 11284 54432
rect 16740 54368 16804 54432
rect 16820 54368 16884 54432
rect 16900 54368 16964 54432
rect 16980 54368 17044 54432
rect 17060 54368 17124 54432
rect 17140 54368 17204 54432
rect 17220 54368 17284 54432
rect 22740 54368 22804 54432
rect 22820 54368 22884 54432
rect 22900 54368 22964 54432
rect 22980 54368 23044 54432
rect 23060 54368 23124 54432
rect 23140 54368 23204 54432
rect 23220 54368 23284 54432
rect 28740 54368 28804 54432
rect 28820 54368 28884 54432
rect 28900 54368 28964 54432
rect 28980 54368 29044 54432
rect 29060 54368 29124 54432
rect 29140 54368 29204 54432
rect 29220 54368 29284 54432
rect 34740 54368 34804 54432
rect 34820 54368 34884 54432
rect 34900 54368 34964 54432
rect 34980 54368 35044 54432
rect 35060 54368 35124 54432
rect 35140 54368 35204 54432
rect 35220 54368 35284 54432
rect 40740 54368 40804 54432
rect 40820 54368 40884 54432
rect 40900 54368 40964 54432
rect 40980 54368 41044 54432
rect 41060 54368 41124 54432
rect 41140 54368 41204 54432
rect 41220 54368 41284 54432
rect 46740 54368 46804 54432
rect 46820 54368 46884 54432
rect 46900 54368 46964 54432
rect 46980 54368 47044 54432
rect 47060 54368 47124 54432
rect 47140 54368 47204 54432
rect 47220 54368 47284 54432
rect 52740 54368 52804 54432
rect 52820 54368 52884 54432
rect 52900 54368 52964 54432
rect 52980 54368 53044 54432
rect 53060 54368 53124 54432
rect 53140 54368 53204 54432
rect 53220 54368 53284 54432
rect 58740 54368 58804 54432
rect 58820 54368 58884 54432
rect 58900 54368 58964 54432
rect 58980 54368 59044 54432
rect 59060 54368 59124 54432
rect 59140 54368 59204 54432
rect 59220 54368 59284 54432
rect 64740 54368 64804 54432
rect 64820 54368 64884 54432
rect 64900 54368 64964 54432
rect 64980 54368 65044 54432
rect 65060 54368 65124 54432
rect 65140 54368 65204 54432
rect 65220 54368 65284 54432
rect 70740 54368 70804 54432
rect 70820 54368 70884 54432
rect 70900 54368 70964 54432
rect 70980 54368 71044 54432
rect 71060 54368 71124 54432
rect 71140 54368 71204 54432
rect 71220 54368 71284 54432
rect 4740 54288 4804 54352
rect 4820 54288 4884 54352
rect 4900 54288 4964 54352
rect 4980 54288 5044 54352
rect 5060 54288 5124 54352
rect 5140 54288 5204 54352
rect 5220 54288 5284 54352
rect 10740 54288 10804 54352
rect 10820 54288 10884 54352
rect 10900 54288 10964 54352
rect 10980 54288 11044 54352
rect 11060 54288 11124 54352
rect 11140 54288 11204 54352
rect 11220 54288 11284 54352
rect 16740 54288 16804 54352
rect 16820 54288 16884 54352
rect 16900 54288 16964 54352
rect 16980 54288 17044 54352
rect 17060 54288 17124 54352
rect 17140 54288 17204 54352
rect 17220 54288 17284 54352
rect 22740 54288 22804 54352
rect 22820 54288 22884 54352
rect 22900 54288 22964 54352
rect 22980 54288 23044 54352
rect 23060 54288 23124 54352
rect 23140 54288 23204 54352
rect 23220 54288 23284 54352
rect 28740 54288 28804 54352
rect 28820 54288 28884 54352
rect 28900 54288 28964 54352
rect 28980 54288 29044 54352
rect 29060 54288 29124 54352
rect 29140 54288 29204 54352
rect 29220 54288 29284 54352
rect 34740 54288 34804 54352
rect 34820 54288 34884 54352
rect 34900 54288 34964 54352
rect 34980 54288 35044 54352
rect 35060 54288 35124 54352
rect 35140 54288 35204 54352
rect 35220 54288 35284 54352
rect 40740 54288 40804 54352
rect 40820 54288 40884 54352
rect 40900 54288 40964 54352
rect 40980 54288 41044 54352
rect 41060 54288 41124 54352
rect 41140 54288 41204 54352
rect 41220 54288 41284 54352
rect 46740 54288 46804 54352
rect 46820 54288 46884 54352
rect 46900 54288 46964 54352
rect 46980 54288 47044 54352
rect 47060 54288 47124 54352
rect 47140 54288 47204 54352
rect 47220 54288 47284 54352
rect 52740 54288 52804 54352
rect 52820 54288 52884 54352
rect 52900 54288 52964 54352
rect 52980 54288 53044 54352
rect 53060 54288 53124 54352
rect 53140 54288 53204 54352
rect 53220 54288 53284 54352
rect 58740 54288 58804 54352
rect 58820 54288 58884 54352
rect 58900 54288 58964 54352
rect 58980 54288 59044 54352
rect 59060 54288 59124 54352
rect 59140 54288 59204 54352
rect 59220 54288 59284 54352
rect 64740 54288 64804 54352
rect 64820 54288 64884 54352
rect 64900 54288 64964 54352
rect 64980 54288 65044 54352
rect 65060 54288 65124 54352
rect 65140 54288 65204 54352
rect 65220 54288 65284 54352
rect 70740 54288 70804 54352
rect 70820 54288 70884 54352
rect 70900 54288 70964 54352
rect 70980 54288 71044 54352
rect 71060 54288 71124 54352
rect 71140 54288 71204 54352
rect 71220 54288 71284 54352
rect 64092 52532 64156 52596
rect 1740 52176 1804 52240
rect 1820 52176 1884 52240
rect 1900 52176 1964 52240
rect 1980 52176 2044 52240
rect 2060 52176 2124 52240
rect 2140 52176 2204 52240
rect 2220 52176 2284 52240
rect 7740 52176 7804 52240
rect 7820 52176 7884 52240
rect 7900 52176 7964 52240
rect 7980 52176 8044 52240
rect 8060 52176 8124 52240
rect 8140 52176 8204 52240
rect 8220 52176 8284 52240
rect 13740 52176 13804 52240
rect 13820 52176 13884 52240
rect 13900 52176 13964 52240
rect 13980 52176 14044 52240
rect 14060 52176 14124 52240
rect 14140 52176 14204 52240
rect 14220 52176 14284 52240
rect 19740 52176 19804 52240
rect 19820 52176 19884 52240
rect 19900 52176 19964 52240
rect 19980 52176 20044 52240
rect 20060 52176 20124 52240
rect 20140 52176 20204 52240
rect 20220 52176 20284 52240
rect 25740 52176 25804 52240
rect 25820 52176 25884 52240
rect 25900 52176 25964 52240
rect 25980 52176 26044 52240
rect 26060 52176 26124 52240
rect 26140 52176 26204 52240
rect 26220 52176 26284 52240
rect 31740 52176 31804 52240
rect 31820 52176 31884 52240
rect 31900 52176 31964 52240
rect 31980 52176 32044 52240
rect 32060 52176 32124 52240
rect 32140 52176 32204 52240
rect 32220 52176 32284 52240
rect 37740 52176 37804 52240
rect 37820 52176 37884 52240
rect 37900 52176 37964 52240
rect 37980 52176 38044 52240
rect 38060 52176 38124 52240
rect 38140 52176 38204 52240
rect 38220 52176 38284 52240
rect 43740 52176 43804 52240
rect 43820 52176 43884 52240
rect 43900 52176 43964 52240
rect 43980 52176 44044 52240
rect 44060 52176 44124 52240
rect 44140 52176 44204 52240
rect 44220 52176 44284 52240
rect 49740 52176 49804 52240
rect 49820 52176 49884 52240
rect 49900 52176 49964 52240
rect 49980 52176 50044 52240
rect 50060 52176 50124 52240
rect 50140 52176 50204 52240
rect 50220 52176 50284 52240
rect 55740 52176 55804 52240
rect 55820 52176 55884 52240
rect 55900 52176 55964 52240
rect 55980 52176 56044 52240
rect 56060 52176 56124 52240
rect 56140 52176 56204 52240
rect 56220 52176 56284 52240
rect 61740 52176 61804 52240
rect 61820 52176 61884 52240
rect 61900 52176 61964 52240
rect 61980 52176 62044 52240
rect 62060 52176 62124 52240
rect 62140 52176 62204 52240
rect 62220 52176 62284 52240
rect 67740 52176 67804 52240
rect 67820 52176 67884 52240
rect 67900 52176 67964 52240
rect 67980 52176 68044 52240
rect 68060 52176 68124 52240
rect 68140 52176 68204 52240
rect 68220 52176 68284 52240
rect 73740 52176 73804 52240
rect 73820 52176 73884 52240
rect 73900 52176 73964 52240
rect 73980 52176 74044 52240
rect 74060 52176 74124 52240
rect 74140 52176 74204 52240
rect 74220 52176 74284 52240
rect 1740 52096 1804 52160
rect 1820 52096 1884 52160
rect 1900 52096 1964 52160
rect 1980 52096 2044 52160
rect 2060 52096 2124 52160
rect 2140 52096 2204 52160
rect 2220 52096 2284 52160
rect 7740 52096 7804 52160
rect 7820 52096 7884 52160
rect 7900 52096 7964 52160
rect 7980 52096 8044 52160
rect 8060 52096 8124 52160
rect 8140 52096 8204 52160
rect 8220 52096 8284 52160
rect 13740 52096 13804 52160
rect 13820 52096 13884 52160
rect 13900 52096 13964 52160
rect 13980 52096 14044 52160
rect 14060 52096 14124 52160
rect 14140 52096 14204 52160
rect 14220 52096 14284 52160
rect 19740 52096 19804 52160
rect 19820 52096 19884 52160
rect 19900 52096 19964 52160
rect 19980 52096 20044 52160
rect 20060 52096 20124 52160
rect 20140 52096 20204 52160
rect 20220 52096 20284 52160
rect 25740 52096 25804 52160
rect 25820 52096 25884 52160
rect 25900 52096 25964 52160
rect 25980 52096 26044 52160
rect 26060 52096 26124 52160
rect 26140 52096 26204 52160
rect 26220 52096 26284 52160
rect 31740 52096 31804 52160
rect 31820 52096 31884 52160
rect 31900 52096 31964 52160
rect 31980 52096 32044 52160
rect 32060 52096 32124 52160
rect 32140 52096 32204 52160
rect 32220 52096 32284 52160
rect 37740 52096 37804 52160
rect 37820 52096 37884 52160
rect 37900 52096 37964 52160
rect 37980 52096 38044 52160
rect 38060 52096 38124 52160
rect 38140 52096 38204 52160
rect 38220 52096 38284 52160
rect 43740 52096 43804 52160
rect 43820 52096 43884 52160
rect 43900 52096 43964 52160
rect 43980 52096 44044 52160
rect 44060 52096 44124 52160
rect 44140 52096 44204 52160
rect 44220 52096 44284 52160
rect 49740 52096 49804 52160
rect 49820 52096 49884 52160
rect 49900 52096 49964 52160
rect 49980 52096 50044 52160
rect 50060 52096 50124 52160
rect 50140 52096 50204 52160
rect 50220 52096 50284 52160
rect 55740 52096 55804 52160
rect 55820 52096 55884 52160
rect 55900 52096 55964 52160
rect 55980 52096 56044 52160
rect 56060 52096 56124 52160
rect 56140 52096 56204 52160
rect 56220 52096 56284 52160
rect 61740 52096 61804 52160
rect 61820 52096 61884 52160
rect 61900 52096 61964 52160
rect 61980 52096 62044 52160
rect 62060 52096 62124 52160
rect 62140 52096 62204 52160
rect 62220 52096 62284 52160
rect 67740 52096 67804 52160
rect 67820 52096 67884 52160
rect 67900 52096 67964 52160
rect 67980 52096 68044 52160
rect 68060 52096 68124 52160
rect 68140 52096 68204 52160
rect 68220 52096 68284 52160
rect 73740 52096 73804 52160
rect 73820 52096 73884 52160
rect 73900 52096 73964 52160
rect 73980 52096 74044 52160
rect 74060 52096 74124 52160
rect 74140 52096 74204 52160
rect 74220 52096 74284 52160
rect 1740 52016 1804 52080
rect 1820 52016 1884 52080
rect 1900 52016 1964 52080
rect 1980 52016 2044 52080
rect 2060 52016 2124 52080
rect 2140 52016 2204 52080
rect 2220 52016 2284 52080
rect 7740 52016 7804 52080
rect 7820 52016 7884 52080
rect 7900 52016 7964 52080
rect 7980 52016 8044 52080
rect 8060 52016 8124 52080
rect 8140 52016 8204 52080
rect 8220 52016 8284 52080
rect 13740 52016 13804 52080
rect 13820 52016 13884 52080
rect 13900 52016 13964 52080
rect 13980 52016 14044 52080
rect 14060 52016 14124 52080
rect 14140 52016 14204 52080
rect 14220 52016 14284 52080
rect 19740 52016 19804 52080
rect 19820 52016 19884 52080
rect 19900 52016 19964 52080
rect 19980 52016 20044 52080
rect 20060 52016 20124 52080
rect 20140 52016 20204 52080
rect 20220 52016 20284 52080
rect 25740 52016 25804 52080
rect 25820 52016 25884 52080
rect 25900 52016 25964 52080
rect 25980 52016 26044 52080
rect 26060 52016 26124 52080
rect 26140 52016 26204 52080
rect 26220 52016 26284 52080
rect 31740 52016 31804 52080
rect 31820 52016 31884 52080
rect 31900 52016 31964 52080
rect 31980 52016 32044 52080
rect 32060 52016 32124 52080
rect 32140 52016 32204 52080
rect 32220 52016 32284 52080
rect 37740 52016 37804 52080
rect 37820 52016 37884 52080
rect 37900 52016 37964 52080
rect 37980 52016 38044 52080
rect 38060 52016 38124 52080
rect 38140 52016 38204 52080
rect 38220 52016 38284 52080
rect 43740 52016 43804 52080
rect 43820 52016 43884 52080
rect 43900 52016 43964 52080
rect 43980 52016 44044 52080
rect 44060 52016 44124 52080
rect 44140 52016 44204 52080
rect 44220 52016 44284 52080
rect 49740 52016 49804 52080
rect 49820 52016 49884 52080
rect 49900 52016 49964 52080
rect 49980 52016 50044 52080
rect 50060 52016 50124 52080
rect 50140 52016 50204 52080
rect 50220 52016 50284 52080
rect 55740 52016 55804 52080
rect 55820 52016 55884 52080
rect 55900 52016 55964 52080
rect 55980 52016 56044 52080
rect 56060 52016 56124 52080
rect 56140 52016 56204 52080
rect 56220 52016 56284 52080
rect 61740 52016 61804 52080
rect 61820 52016 61884 52080
rect 61900 52016 61964 52080
rect 61980 52016 62044 52080
rect 62060 52016 62124 52080
rect 62140 52016 62204 52080
rect 62220 52016 62284 52080
rect 67740 52016 67804 52080
rect 67820 52016 67884 52080
rect 67900 52016 67964 52080
rect 67980 52016 68044 52080
rect 68060 52016 68124 52080
rect 68140 52016 68204 52080
rect 68220 52016 68284 52080
rect 73740 52016 73804 52080
rect 73820 52016 73884 52080
rect 73900 52016 73964 52080
rect 73980 52016 74044 52080
rect 74060 52016 74124 52080
rect 74140 52016 74204 52080
rect 74220 52016 74284 52080
rect 1740 51936 1804 52000
rect 1820 51936 1884 52000
rect 1900 51936 1964 52000
rect 1980 51936 2044 52000
rect 2060 51936 2124 52000
rect 2140 51936 2204 52000
rect 2220 51936 2284 52000
rect 7740 51936 7804 52000
rect 7820 51936 7884 52000
rect 7900 51936 7964 52000
rect 7980 51936 8044 52000
rect 8060 51936 8124 52000
rect 8140 51936 8204 52000
rect 8220 51936 8284 52000
rect 13740 51936 13804 52000
rect 13820 51936 13884 52000
rect 13900 51936 13964 52000
rect 13980 51936 14044 52000
rect 14060 51936 14124 52000
rect 14140 51936 14204 52000
rect 14220 51936 14284 52000
rect 19740 51936 19804 52000
rect 19820 51936 19884 52000
rect 19900 51936 19964 52000
rect 19980 51936 20044 52000
rect 20060 51936 20124 52000
rect 20140 51936 20204 52000
rect 20220 51936 20284 52000
rect 25740 51936 25804 52000
rect 25820 51936 25884 52000
rect 25900 51936 25964 52000
rect 25980 51936 26044 52000
rect 26060 51936 26124 52000
rect 26140 51936 26204 52000
rect 26220 51936 26284 52000
rect 31740 51936 31804 52000
rect 31820 51936 31884 52000
rect 31900 51936 31964 52000
rect 31980 51936 32044 52000
rect 32060 51936 32124 52000
rect 32140 51936 32204 52000
rect 32220 51936 32284 52000
rect 37740 51936 37804 52000
rect 37820 51936 37884 52000
rect 37900 51936 37964 52000
rect 37980 51936 38044 52000
rect 38060 51936 38124 52000
rect 38140 51936 38204 52000
rect 38220 51936 38284 52000
rect 43740 51936 43804 52000
rect 43820 51936 43884 52000
rect 43900 51936 43964 52000
rect 43980 51936 44044 52000
rect 44060 51936 44124 52000
rect 44140 51936 44204 52000
rect 44220 51936 44284 52000
rect 49740 51936 49804 52000
rect 49820 51936 49884 52000
rect 49900 51936 49964 52000
rect 49980 51936 50044 52000
rect 50060 51936 50124 52000
rect 50140 51936 50204 52000
rect 50220 51936 50284 52000
rect 55740 51936 55804 52000
rect 55820 51936 55884 52000
rect 55900 51936 55964 52000
rect 55980 51936 56044 52000
rect 56060 51936 56124 52000
rect 56140 51936 56204 52000
rect 56220 51936 56284 52000
rect 61740 51936 61804 52000
rect 61820 51936 61884 52000
rect 61900 51936 61964 52000
rect 61980 51936 62044 52000
rect 62060 51936 62124 52000
rect 62140 51936 62204 52000
rect 62220 51936 62284 52000
rect 67740 51936 67804 52000
rect 67820 51936 67884 52000
rect 67900 51936 67964 52000
rect 67980 51936 68044 52000
rect 68060 51936 68124 52000
rect 68140 51936 68204 52000
rect 68220 51936 68284 52000
rect 73740 51936 73804 52000
rect 73820 51936 73884 52000
rect 73900 51936 73964 52000
rect 73980 51936 74044 52000
rect 74060 51936 74124 52000
rect 74140 51936 74204 52000
rect 74220 51936 74284 52000
rect 64276 50220 64340 50284
rect 62988 48724 63052 48788
rect 64460 48044 64524 48108
rect 63908 47696 63972 47700
rect 63908 47640 63922 47696
rect 63922 47640 63972 47696
rect 63908 47636 63972 47640
rect 4740 44528 4804 44592
rect 4820 44528 4884 44592
rect 4900 44528 4964 44592
rect 4980 44528 5044 44592
rect 5060 44528 5124 44592
rect 5140 44528 5204 44592
rect 5220 44528 5284 44592
rect 10740 44528 10804 44592
rect 10820 44528 10884 44592
rect 10900 44528 10964 44592
rect 10980 44528 11044 44592
rect 11060 44528 11124 44592
rect 11140 44528 11204 44592
rect 11220 44528 11284 44592
rect 16740 44528 16804 44592
rect 16820 44528 16884 44592
rect 16900 44528 16964 44592
rect 16980 44528 17044 44592
rect 17060 44528 17124 44592
rect 17140 44528 17204 44592
rect 17220 44528 17284 44592
rect 22740 44528 22804 44592
rect 22820 44528 22884 44592
rect 22900 44528 22964 44592
rect 22980 44528 23044 44592
rect 23060 44528 23124 44592
rect 23140 44528 23204 44592
rect 23220 44528 23284 44592
rect 28740 44528 28804 44592
rect 28820 44528 28884 44592
rect 28900 44528 28964 44592
rect 28980 44528 29044 44592
rect 29060 44528 29124 44592
rect 29140 44528 29204 44592
rect 29220 44528 29284 44592
rect 34740 44528 34804 44592
rect 34820 44528 34884 44592
rect 34900 44528 34964 44592
rect 34980 44528 35044 44592
rect 35060 44528 35124 44592
rect 35140 44528 35204 44592
rect 35220 44528 35284 44592
rect 40740 44528 40804 44592
rect 40820 44528 40884 44592
rect 40900 44528 40964 44592
rect 40980 44528 41044 44592
rect 41060 44528 41124 44592
rect 41140 44528 41204 44592
rect 41220 44528 41284 44592
rect 46740 44528 46804 44592
rect 46820 44528 46884 44592
rect 46900 44528 46964 44592
rect 46980 44528 47044 44592
rect 47060 44528 47124 44592
rect 47140 44528 47204 44592
rect 47220 44528 47284 44592
rect 52740 44528 52804 44592
rect 52820 44528 52884 44592
rect 52900 44528 52964 44592
rect 52980 44528 53044 44592
rect 53060 44528 53124 44592
rect 53140 44528 53204 44592
rect 53220 44528 53284 44592
rect 58740 44528 58804 44592
rect 58820 44528 58884 44592
rect 58900 44528 58964 44592
rect 58980 44528 59044 44592
rect 59060 44528 59124 44592
rect 59140 44528 59204 44592
rect 59220 44528 59284 44592
rect 64740 44528 64804 44592
rect 64820 44528 64884 44592
rect 64900 44528 64964 44592
rect 64980 44528 65044 44592
rect 65060 44528 65124 44592
rect 65140 44528 65204 44592
rect 65220 44528 65284 44592
rect 70740 44528 70804 44592
rect 70820 44528 70884 44592
rect 70900 44528 70964 44592
rect 70980 44528 71044 44592
rect 71060 44528 71124 44592
rect 71140 44528 71204 44592
rect 71220 44528 71284 44592
rect 4740 44448 4804 44512
rect 4820 44448 4884 44512
rect 4900 44448 4964 44512
rect 4980 44448 5044 44512
rect 5060 44448 5124 44512
rect 5140 44448 5204 44512
rect 5220 44448 5284 44512
rect 10740 44448 10804 44512
rect 10820 44448 10884 44512
rect 10900 44448 10964 44512
rect 10980 44448 11044 44512
rect 11060 44448 11124 44512
rect 11140 44448 11204 44512
rect 11220 44448 11284 44512
rect 16740 44448 16804 44512
rect 16820 44448 16884 44512
rect 16900 44448 16964 44512
rect 16980 44448 17044 44512
rect 17060 44448 17124 44512
rect 17140 44448 17204 44512
rect 17220 44448 17284 44512
rect 22740 44448 22804 44512
rect 22820 44448 22884 44512
rect 22900 44448 22964 44512
rect 22980 44448 23044 44512
rect 23060 44448 23124 44512
rect 23140 44448 23204 44512
rect 23220 44448 23284 44512
rect 28740 44448 28804 44512
rect 28820 44448 28884 44512
rect 28900 44448 28964 44512
rect 28980 44448 29044 44512
rect 29060 44448 29124 44512
rect 29140 44448 29204 44512
rect 29220 44448 29284 44512
rect 34740 44448 34804 44512
rect 34820 44448 34884 44512
rect 34900 44448 34964 44512
rect 34980 44448 35044 44512
rect 35060 44448 35124 44512
rect 35140 44448 35204 44512
rect 35220 44448 35284 44512
rect 40740 44448 40804 44512
rect 40820 44448 40884 44512
rect 40900 44448 40964 44512
rect 40980 44448 41044 44512
rect 41060 44448 41124 44512
rect 41140 44448 41204 44512
rect 41220 44448 41284 44512
rect 46740 44448 46804 44512
rect 46820 44448 46884 44512
rect 46900 44448 46964 44512
rect 46980 44448 47044 44512
rect 47060 44448 47124 44512
rect 47140 44448 47204 44512
rect 47220 44448 47284 44512
rect 52740 44448 52804 44512
rect 52820 44448 52884 44512
rect 52900 44448 52964 44512
rect 52980 44448 53044 44512
rect 53060 44448 53124 44512
rect 53140 44448 53204 44512
rect 53220 44448 53284 44512
rect 58740 44448 58804 44512
rect 58820 44448 58884 44512
rect 58900 44448 58964 44512
rect 58980 44448 59044 44512
rect 59060 44448 59124 44512
rect 59140 44448 59204 44512
rect 59220 44448 59284 44512
rect 64740 44448 64804 44512
rect 64820 44448 64884 44512
rect 64900 44448 64964 44512
rect 64980 44448 65044 44512
rect 65060 44448 65124 44512
rect 65140 44448 65204 44512
rect 65220 44448 65284 44512
rect 70740 44448 70804 44512
rect 70820 44448 70884 44512
rect 70900 44448 70964 44512
rect 70980 44448 71044 44512
rect 71060 44448 71124 44512
rect 71140 44448 71204 44512
rect 71220 44448 71284 44512
rect 4740 44368 4804 44432
rect 4820 44368 4884 44432
rect 4900 44368 4964 44432
rect 4980 44368 5044 44432
rect 5060 44368 5124 44432
rect 5140 44368 5204 44432
rect 5220 44368 5284 44432
rect 10740 44368 10804 44432
rect 10820 44368 10884 44432
rect 10900 44368 10964 44432
rect 10980 44368 11044 44432
rect 11060 44368 11124 44432
rect 11140 44368 11204 44432
rect 11220 44368 11284 44432
rect 16740 44368 16804 44432
rect 16820 44368 16884 44432
rect 16900 44368 16964 44432
rect 16980 44368 17044 44432
rect 17060 44368 17124 44432
rect 17140 44368 17204 44432
rect 17220 44368 17284 44432
rect 22740 44368 22804 44432
rect 22820 44368 22884 44432
rect 22900 44368 22964 44432
rect 22980 44368 23044 44432
rect 23060 44368 23124 44432
rect 23140 44368 23204 44432
rect 23220 44368 23284 44432
rect 28740 44368 28804 44432
rect 28820 44368 28884 44432
rect 28900 44368 28964 44432
rect 28980 44368 29044 44432
rect 29060 44368 29124 44432
rect 29140 44368 29204 44432
rect 29220 44368 29284 44432
rect 34740 44368 34804 44432
rect 34820 44368 34884 44432
rect 34900 44368 34964 44432
rect 34980 44368 35044 44432
rect 35060 44368 35124 44432
rect 35140 44368 35204 44432
rect 35220 44368 35284 44432
rect 40740 44368 40804 44432
rect 40820 44368 40884 44432
rect 40900 44368 40964 44432
rect 40980 44368 41044 44432
rect 41060 44368 41124 44432
rect 41140 44368 41204 44432
rect 41220 44368 41284 44432
rect 46740 44368 46804 44432
rect 46820 44368 46884 44432
rect 46900 44368 46964 44432
rect 46980 44368 47044 44432
rect 47060 44368 47124 44432
rect 47140 44368 47204 44432
rect 47220 44368 47284 44432
rect 52740 44368 52804 44432
rect 52820 44368 52884 44432
rect 52900 44368 52964 44432
rect 52980 44368 53044 44432
rect 53060 44368 53124 44432
rect 53140 44368 53204 44432
rect 53220 44368 53284 44432
rect 58740 44368 58804 44432
rect 58820 44368 58884 44432
rect 58900 44368 58964 44432
rect 58980 44368 59044 44432
rect 59060 44368 59124 44432
rect 59140 44368 59204 44432
rect 59220 44368 59284 44432
rect 64740 44368 64804 44432
rect 64820 44368 64884 44432
rect 64900 44368 64964 44432
rect 64980 44368 65044 44432
rect 65060 44368 65124 44432
rect 65140 44368 65204 44432
rect 65220 44368 65284 44432
rect 70740 44368 70804 44432
rect 70820 44368 70884 44432
rect 70900 44368 70964 44432
rect 70980 44368 71044 44432
rect 71060 44368 71124 44432
rect 71140 44368 71204 44432
rect 71220 44368 71284 44432
rect 4740 44288 4804 44352
rect 4820 44288 4884 44352
rect 4900 44288 4964 44352
rect 4980 44288 5044 44352
rect 5060 44288 5124 44352
rect 5140 44288 5204 44352
rect 5220 44288 5284 44352
rect 10740 44288 10804 44352
rect 10820 44288 10884 44352
rect 10900 44288 10964 44352
rect 10980 44288 11044 44352
rect 11060 44288 11124 44352
rect 11140 44288 11204 44352
rect 11220 44288 11284 44352
rect 16740 44288 16804 44352
rect 16820 44288 16884 44352
rect 16900 44288 16964 44352
rect 16980 44288 17044 44352
rect 17060 44288 17124 44352
rect 17140 44288 17204 44352
rect 17220 44288 17284 44352
rect 22740 44288 22804 44352
rect 22820 44288 22884 44352
rect 22900 44288 22964 44352
rect 22980 44288 23044 44352
rect 23060 44288 23124 44352
rect 23140 44288 23204 44352
rect 23220 44288 23284 44352
rect 28740 44288 28804 44352
rect 28820 44288 28884 44352
rect 28900 44288 28964 44352
rect 28980 44288 29044 44352
rect 29060 44288 29124 44352
rect 29140 44288 29204 44352
rect 29220 44288 29284 44352
rect 34740 44288 34804 44352
rect 34820 44288 34884 44352
rect 34900 44288 34964 44352
rect 34980 44288 35044 44352
rect 35060 44288 35124 44352
rect 35140 44288 35204 44352
rect 35220 44288 35284 44352
rect 40740 44288 40804 44352
rect 40820 44288 40884 44352
rect 40900 44288 40964 44352
rect 40980 44288 41044 44352
rect 41060 44288 41124 44352
rect 41140 44288 41204 44352
rect 41220 44288 41284 44352
rect 46740 44288 46804 44352
rect 46820 44288 46884 44352
rect 46900 44288 46964 44352
rect 46980 44288 47044 44352
rect 47060 44288 47124 44352
rect 47140 44288 47204 44352
rect 47220 44288 47284 44352
rect 52740 44288 52804 44352
rect 52820 44288 52884 44352
rect 52900 44288 52964 44352
rect 52980 44288 53044 44352
rect 53060 44288 53124 44352
rect 53140 44288 53204 44352
rect 53220 44288 53284 44352
rect 58740 44288 58804 44352
rect 58820 44288 58884 44352
rect 58900 44288 58964 44352
rect 58980 44288 59044 44352
rect 59060 44288 59124 44352
rect 59140 44288 59204 44352
rect 59220 44288 59284 44352
rect 64740 44288 64804 44352
rect 64820 44288 64884 44352
rect 64900 44288 64964 44352
rect 64980 44288 65044 44352
rect 65060 44288 65124 44352
rect 65140 44288 65204 44352
rect 65220 44288 65284 44352
rect 70740 44288 70804 44352
rect 70820 44288 70884 44352
rect 70900 44288 70964 44352
rect 70980 44288 71044 44352
rect 71060 44288 71124 44352
rect 71140 44288 71204 44352
rect 71220 44288 71284 44352
rect 1740 42176 1804 42240
rect 1820 42176 1884 42240
rect 1900 42176 1964 42240
rect 1980 42176 2044 42240
rect 2060 42176 2124 42240
rect 2140 42176 2204 42240
rect 2220 42176 2284 42240
rect 7740 42176 7804 42240
rect 7820 42176 7884 42240
rect 7900 42176 7964 42240
rect 7980 42176 8044 42240
rect 8060 42176 8124 42240
rect 8140 42176 8204 42240
rect 8220 42176 8284 42240
rect 13740 42176 13804 42240
rect 13820 42176 13884 42240
rect 13900 42176 13964 42240
rect 13980 42176 14044 42240
rect 14060 42176 14124 42240
rect 14140 42176 14204 42240
rect 14220 42176 14284 42240
rect 19740 42176 19804 42240
rect 19820 42176 19884 42240
rect 19900 42176 19964 42240
rect 19980 42176 20044 42240
rect 20060 42176 20124 42240
rect 20140 42176 20204 42240
rect 20220 42176 20284 42240
rect 25740 42176 25804 42240
rect 25820 42176 25884 42240
rect 25900 42176 25964 42240
rect 25980 42176 26044 42240
rect 26060 42176 26124 42240
rect 26140 42176 26204 42240
rect 26220 42176 26284 42240
rect 31740 42176 31804 42240
rect 31820 42176 31884 42240
rect 31900 42176 31964 42240
rect 31980 42176 32044 42240
rect 32060 42176 32124 42240
rect 32140 42176 32204 42240
rect 32220 42176 32284 42240
rect 37740 42176 37804 42240
rect 37820 42176 37884 42240
rect 37900 42176 37964 42240
rect 37980 42176 38044 42240
rect 38060 42176 38124 42240
rect 38140 42176 38204 42240
rect 38220 42176 38284 42240
rect 43740 42176 43804 42240
rect 43820 42176 43884 42240
rect 43900 42176 43964 42240
rect 43980 42176 44044 42240
rect 44060 42176 44124 42240
rect 44140 42176 44204 42240
rect 44220 42176 44284 42240
rect 49740 42176 49804 42240
rect 49820 42176 49884 42240
rect 49900 42176 49964 42240
rect 49980 42176 50044 42240
rect 50060 42176 50124 42240
rect 50140 42176 50204 42240
rect 50220 42176 50284 42240
rect 55740 42176 55804 42240
rect 55820 42176 55884 42240
rect 55900 42176 55964 42240
rect 55980 42176 56044 42240
rect 56060 42176 56124 42240
rect 56140 42176 56204 42240
rect 56220 42176 56284 42240
rect 61740 42176 61804 42240
rect 61820 42176 61884 42240
rect 61900 42176 61964 42240
rect 61980 42176 62044 42240
rect 62060 42176 62124 42240
rect 62140 42176 62204 42240
rect 62220 42176 62284 42240
rect 67740 42176 67804 42240
rect 67820 42176 67884 42240
rect 67900 42176 67964 42240
rect 67980 42176 68044 42240
rect 68060 42176 68124 42240
rect 68140 42176 68204 42240
rect 68220 42176 68284 42240
rect 73740 42176 73804 42240
rect 73820 42176 73884 42240
rect 73900 42176 73964 42240
rect 73980 42176 74044 42240
rect 74060 42176 74124 42240
rect 74140 42176 74204 42240
rect 74220 42176 74284 42240
rect 1740 42096 1804 42160
rect 1820 42096 1884 42160
rect 1900 42096 1964 42160
rect 1980 42096 2044 42160
rect 2060 42096 2124 42160
rect 2140 42096 2204 42160
rect 2220 42096 2284 42160
rect 7740 42096 7804 42160
rect 7820 42096 7884 42160
rect 7900 42096 7964 42160
rect 7980 42096 8044 42160
rect 8060 42096 8124 42160
rect 8140 42096 8204 42160
rect 8220 42096 8284 42160
rect 13740 42096 13804 42160
rect 13820 42096 13884 42160
rect 13900 42096 13964 42160
rect 13980 42096 14044 42160
rect 14060 42096 14124 42160
rect 14140 42096 14204 42160
rect 14220 42096 14284 42160
rect 19740 42096 19804 42160
rect 19820 42096 19884 42160
rect 19900 42096 19964 42160
rect 19980 42096 20044 42160
rect 20060 42096 20124 42160
rect 20140 42096 20204 42160
rect 20220 42096 20284 42160
rect 25740 42096 25804 42160
rect 25820 42096 25884 42160
rect 25900 42096 25964 42160
rect 25980 42096 26044 42160
rect 26060 42096 26124 42160
rect 26140 42096 26204 42160
rect 26220 42096 26284 42160
rect 31740 42096 31804 42160
rect 31820 42096 31884 42160
rect 31900 42096 31964 42160
rect 31980 42096 32044 42160
rect 32060 42096 32124 42160
rect 32140 42096 32204 42160
rect 32220 42096 32284 42160
rect 37740 42096 37804 42160
rect 37820 42096 37884 42160
rect 37900 42096 37964 42160
rect 37980 42096 38044 42160
rect 38060 42096 38124 42160
rect 38140 42096 38204 42160
rect 38220 42096 38284 42160
rect 43740 42096 43804 42160
rect 43820 42096 43884 42160
rect 43900 42096 43964 42160
rect 43980 42096 44044 42160
rect 44060 42096 44124 42160
rect 44140 42096 44204 42160
rect 44220 42096 44284 42160
rect 49740 42096 49804 42160
rect 49820 42096 49884 42160
rect 49900 42096 49964 42160
rect 49980 42096 50044 42160
rect 50060 42096 50124 42160
rect 50140 42096 50204 42160
rect 50220 42096 50284 42160
rect 55740 42096 55804 42160
rect 55820 42096 55884 42160
rect 55900 42096 55964 42160
rect 55980 42096 56044 42160
rect 56060 42096 56124 42160
rect 56140 42096 56204 42160
rect 56220 42096 56284 42160
rect 61740 42096 61804 42160
rect 61820 42096 61884 42160
rect 61900 42096 61964 42160
rect 61980 42096 62044 42160
rect 62060 42096 62124 42160
rect 62140 42096 62204 42160
rect 62220 42096 62284 42160
rect 67740 42096 67804 42160
rect 67820 42096 67884 42160
rect 67900 42096 67964 42160
rect 67980 42096 68044 42160
rect 68060 42096 68124 42160
rect 68140 42096 68204 42160
rect 68220 42096 68284 42160
rect 73740 42096 73804 42160
rect 73820 42096 73884 42160
rect 73900 42096 73964 42160
rect 73980 42096 74044 42160
rect 74060 42096 74124 42160
rect 74140 42096 74204 42160
rect 74220 42096 74284 42160
rect 1740 42016 1804 42080
rect 1820 42016 1884 42080
rect 1900 42016 1964 42080
rect 1980 42016 2044 42080
rect 2060 42016 2124 42080
rect 2140 42016 2204 42080
rect 2220 42016 2284 42080
rect 7740 42016 7804 42080
rect 7820 42016 7884 42080
rect 7900 42016 7964 42080
rect 7980 42016 8044 42080
rect 8060 42016 8124 42080
rect 8140 42016 8204 42080
rect 8220 42016 8284 42080
rect 13740 42016 13804 42080
rect 13820 42016 13884 42080
rect 13900 42016 13964 42080
rect 13980 42016 14044 42080
rect 14060 42016 14124 42080
rect 14140 42016 14204 42080
rect 14220 42016 14284 42080
rect 19740 42016 19804 42080
rect 19820 42016 19884 42080
rect 19900 42016 19964 42080
rect 19980 42016 20044 42080
rect 20060 42016 20124 42080
rect 20140 42016 20204 42080
rect 20220 42016 20284 42080
rect 25740 42016 25804 42080
rect 25820 42016 25884 42080
rect 25900 42016 25964 42080
rect 25980 42016 26044 42080
rect 26060 42016 26124 42080
rect 26140 42016 26204 42080
rect 26220 42016 26284 42080
rect 31740 42016 31804 42080
rect 31820 42016 31884 42080
rect 31900 42016 31964 42080
rect 31980 42016 32044 42080
rect 32060 42016 32124 42080
rect 32140 42016 32204 42080
rect 32220 42016 32284 42080
rect 37740 42016 37804 42080
rect 37820 42016 37884 42080
rect 37900 42016 37964 42080
rect 37980 42016 38044 42080
rect 38060 42016 38124 42080
rect 38140 42016 38204 42080
rect 38220 42016 38284 42080
rect 43740 42016 43804 42080
rect 43820 42016 43884 42080
rect 43900 42016 43964 42080
rect 43980 42016 44044 42080
rect 44060 42016 44124 42080
rect 44140 42016 44204 42080
rect 44220 42016 44284 42080
rect 49740 42016 49804 42080
rect 49820 42016 49884 42080
rect 49900 42016 49964 42080
rect 49980 42016 50044 42080
rect 50060 42016 50124 42080
rect 50140 42016 50204 42080
rect 50220 42016 50284 42080
rect 55740 42016 55804 42080
rect 55820 42016 55884 42080
rect 55900 42016 55964 42080
rect 55980 42016 56044 42080
rect 56060 42016 56124 42080
rect 56140 42016 56204 42080
rect 56220 42016 56284 42080
rect 61740 42016 61804 42080
rect 61820 42016 61884 42080
rect 61900 42016 61964 42080
rect 61980 42016 62044 42080
rect 62060 42016 62124 42080
rect 62140 42016 62204 42080
rect 62220 42016 62284 42080
rect 67740 42016 67804 42080
rect 67820 42016 67884 42080
rect 67900 42016 67964 42080
rect 67980 42016 68044 42080
rect 68060 42016 68124 42080
rect 68140 42016 68204 42080
rect 68220 42016 68284 42080
rect 73740 42016 73804 42080
rect 73820 42016 73884 42080
rect 73900 42016 73964 42080
rect 73980 42016 74044 42080
rect 74060 42016 74124 42080
rect 74140 42016 74204 42080
rect 74220 42016 74284 42080
rect 1740 41936 1804 42000
rect 1820 41936 1884 42000
rect 1900 41936 1964 42000
rect 1980 41936 2044 42000
rect 2060 41936 2124 42000
rect 2140 41936 2204 42000
rect 2220 41936 2284 42000
rect 7740 41936 7804 42000
rect 7820 41936 7884 42000
rect 7900 41936 7964 42000
rect 7980 41936 8044 42000
rect 8060 41936 8124 42000
rect 8140 41936 8204 42000
rect 8220 41936 8284 42000
rect 13740 41936 13804 42000
rect 13820 41936 13884 42000
rect 13900 41936 13964 42000
rect 13980 41936 14044 42000
rect 14060 41936 14124 42000
rect 14140 41936 14204 42000
rect 14220 41936 14284 42000
rect 19740 41936 19804 42000
rect 19820 41936 19884 42000
rect 19900 41936 19964 42000
rect 19980 41936 20044 42000
rect 20060 41936 20124 42000
rect 20140 41936 20204 42000
rect 20220 41936 20284 42000
rect 25740 41936 25804 42000
rect 25820 41936 25884 42000
rect 25900 41936 25964 42000
rect 25980 41936 26044 42000
rect 26060 41936 26124 42000
rect 26140 41936 26204 42000
rect 26220 41936 26284 42000
rect 31740 41936 31804 42000
rect 31820 41936 31884 42000
rect 31900 41936 31964 42000
rect 31980 41936 32044 42000
rect 32060 41936 32124 42000
rect 32140 41936 32204 42000
rect 32220 41936 32284 42000
rect 37740 41936 37804 42000
rect 37820 41936 37884 42000
rect 37900 41936 37964 42000
rect 37980 41936 38044 42000
rect 38060 41936 38124 42000
rect 38140 41936 38204 42000
rect 38220 41936 38284 42000
rect 43740 41936 43804 42000
rect 43820 41936 43884 42000
rect 43900 41936 43964 42000
rect 43980 41936 44044 42000
rect 44060 41936 44124 42000
rect 44140 41936 44204 42000
rect 44220 41936 44284 42000
rect 49740 41936 49804 42000
rect 49820 41936 49884 42000
rect 49900 41936 49964 42000
rect 49980 41936 50044 42000
rect 50060 41936 50124 42000
rect 50140 41936 50204 42000
rect 50220 41936 50284 42000
rect 55740 41936 55804 42000
rect 55820 41936 55884 42000
rect 55900 41936 55964 42000
rect 55980 41936 56044 42000
rect 56060 41936 56124 42000
rect 56140 41936 56204 42000
rect 56220 41936 56284 42000
rect 61740 41936 61804 42000
rect 61820 41936 61884 42000
rect 61900 41936 61964 42000
rect 61980 41936 62044 42000
rect 62060 41936 62124 42000
rect 62140 41936 62204 42000
rect 62220 41936 62284 42000
rect 67740 41936 67804 42000
rect 67820 41936 67884 42000
rect 67900 41936 67964 42000
rect 67980 41936 68044 42000
rect 68060 41936 68124 42000
rect 68140 41936 68204 42000
rect 68220 41936 68284 42000
rect 73740 41936 73804 42000
rect 73820 41936 73884 42000
rect 73900 41936 73964 42000
rect 73980 41936 74044 42000
rect 74060 41936 74124 42000
rect 74140 41936 74204 42000
rect 74220 41936 74284 42000
rect 65564 40836 65628 40900
rect 65748 38796 65812 38860
rect 65932 34716 65996 34780
rect 4740 34528 4804 34592
rect 4820 34528 4884 34592
rect 4900 34528 4964 34592
rect 4980 34528 5044 34592
rect 5060 34528 5124 34592
rect 5140 34528 5204 34592
rect 5220 34528 5284 34592
rect 10740 34528 10804 34592
rect 10820 34528 10884 34592
rect 10900 34528 10964 34592
rect 10980 34528 11044 34592
rect 11060 34528 11124 34592
rect 11140 34528 11204 34592
rect 11220 34528 11284 34592
rect 16740 34528 16804 34592
rect 16820 34528 16884 34592
rect 16900 34528 16964 34592
rect 16980 34528 17044 34592
rect 17060 34528 17124 34592
rect 17140 34528 17204 34592
rect 17220 34528 17284 34592
rect 22740 34528 22804 34592
rect 22820 34528 22884 34592
rect 22900 34528 22964 34592
rect 22980 34528 23044 34592
rect 23060 34528 23124 34592
rect 23140 34528 23204 34592
rect 23220 34528 23284 34592
rect 28740 34528 28804 34592
rect 28820 34528 28884 34592
rect 28900 34528 28964 34592
rect 28980 34528 29044 34592
rect 29060 34528 29124 34592
rect 29140 34528 29204 34592
rect 29220 34528 29284 34592
rect 34740 34528 34804 34592
rect 34820 34528 34884 34592
rect 34900 34528 34964 34592
rect 34980 34528 35044 34592
rect 35060 34528 35124 34592
rect 35140 34528 35204 34592
rect 35220 34528 35284 34592
rect 40740 34528 40804 34592
rect 40820 34528 40884 34592
rect 40900 34528 40964 34592
rect 40980 34528 41044 34592
rect 41060 34528 41124 34592
rect 41140 34528 41204 34592
rect 41220 34528 41284 34592
rect 46740 34528 46804 34592
rect 46820 34528 46884 34592
rect 46900 34528 46964 34592
rect 46980 34528 47044 34592
rect 47060 34528 47124 34592
rect 47140 34528 47204 34592
rect 47220 34528 47284 34592
rect 52740 34528 52804 34592
rect 52820 34528 52884 34592
rect 52900 34528 52964 34592
rect 52980 34528 53044 34592
rect 53060 34528 53124 34592
rect 53140 34528 53204 34592
rect 53220 34528 53284 34592
rect 58740 34528 58804 34592
rect 58820 34528 58884 34592
rect 58900 34528 58964 34592
rect 58980 34528 59044 34592
rect 59060 34528 59124 34592
rect 59140 34528 59204 34592
rect 59220 34528 59284 34592
rect 64740 34528 64804 34592
rect 64820 34528 64884 34592
rect 64900 34528 64964 34592
rect 64980 34528 65044 34592
rect 65060 34528 65124 34592
rect 65140 34528 65204 34592
rect 65220 34528 65284 34592
rect 70740 34528 70804 34592
rect 70820 34528 70884 34592
rect 70900 34528 70964 34592
rect 70980 34528 71044 34592
rect 71060 34528 71124 34592
rect 71140 34528 71204 34592
rect 71220 34528 71284 34592
rect 4740 34448 4804 34512
rect 4820 34448 4884 34512
rect 4900 34448 4964 34512
rect 4980 34448 5044 34512
rect 5060 34448 5124 34512
rect 5140 34448 5204 34512
rect 5220 34448 5284 34512
rect 10740 34448 10804 34512
rect 10820 34448 10884 34512
rect 10900 34448 10964 34512
rect 10980 34448 11044 34512
rect 11060 34448 11124 34512
rect 11140 34448 11204 34512
rect 11220 34448 11284 34512
rect 16740 34448 16804 34512
rect 16820 34448 16884 34512
rect 16900 34448 16964 34512
rect 16980 34448 17044 34512
rect 17060 34448 17124 34512
rect 17140 34448 17204 34512
rect 17220 34448 17284 34512
rect 22740 34448 22804 34512
rect 22820 34448 22884 34512
rect 22900 34448 22964 34512
rect 22980 34448 23044 34512
rect 23060 34448 23124 34512
rect 23140 34448 23204 34512
rect 23220 34448 23284 34512
rect 28740 34448 28804 34512
rect 28820 34448 28884 34512
rect 28900 34448 28964 34512
rect 28980 34448 29044 34512
rect 29060 34448 29124 34512
rect 29140 34448 29204 34512
rect 29220 34448 29284 34512
rect 34740 34448 34804 34512
rect 34820 34448 34884 34512
rect 34900 34448 34964 34512
rect 34980 34448 35044 34512
rect 35060 34448 35124 34512
rect 35140 34448 35204 34512
rect 35220 34448 35284 34512
rect 40740 34448 40804 34512
rect 40820 34448 40884 34512
rect 40900 34448 40964 34512
rect 40980 34448 41044 34512
rect 41060 34448 41124 34512
rect 41140 34448 41204 34512
rect 41220 34448 41284 34512
rect 46740 34448 46804 34512
rect 46820 34448 46884 34512
rect 46900 34448 46964 34512
rect 46980 34448 47044 34512
rect 47060 34448 47124 34512
rect 47140 34448 47204 34512
rect 47220 34448 47284 34512
rect 52740 34448 52804 34512
rect 52820 34448 52884 34512
rect 52900 34448 52964 34512
rect 52980 34448 53044 34512
rect 53060 34448 53124 34512
rect 53140 34448 53204 34512
rect 53220 34448 53284 34512
rect 58740 34448 58804 34512
rect 58820 34448 58884 34512
rect 58900 34448 58964 34512
rect 58980 34448 59044 34512
rect 59060 34448 59124 34512
rect 59140 34448 59204 34512
rect 59220 34448 59284 34512
rect 64740 34448 64804 34512
rect 64820 34448 64884 34512
rect 64900 34448 64964 34512
rect 64980 34448 65044 34512
rect 65060 34448 65124 34512
rect 65140 34448 65204 34512
rect 65220 34448 65284 34512
rect 70740 34448 70804 34512
rect 70820 34448 70884 34512
rect 70900 34448 70964 34512
rect 70980 34448 71044 34512
rect 71060 34448 71124 34512
rect 71140 34448 71204 34512
rect 71220 34448 71284 34512
rect 4740 34368 4804 34432
rect 4820 34368 4884 34432
rect 4900 34368 4964 34432
rect 4980 34368 5044 34432
rect 5060 34368 5124 34432
rect 5140 34368 5204 34432
rect 5220 34368 5284 34432
rect 10740 34368 10804 34432
rect 10820 34368 10884 34432
rect 10900 34368 10964 34432
rect 10980 34368 11044 34432
rect 11060 34368 11124 34432
rect 11140 34368 11204 34432
rect 11220 34368 11284 34432
rect 16740 34368 16804 34432
rect 16820 34368 16884 34432
rect 16900 34368 16964 34432
rect 16980 34368 17044 34432
rect 17060 34368 17124 34432
rect 17140 34368 17204 34432
rect 17220 34368 17284 34432
rect 22740 34368 22804 34432
rect 22820 34368 22884 34432
rect 22900 34368 22964 34432
rect 22980 34368 23044 34432
rect 23060 34368 23124 34432
rect 23140 34368 23204 34432
rect 23220 34368 23284 34432
rect 28740 34368 28804 34432
rect 28820 34368 28884 34432
rect 28900 34368 28964 34432
rect 28980 34368 29044 34432
rect 29060 34368 29124 34432
rect 29140 34368 29204 34432
rect 29220 34368 29284 34432
rect 34740 34368 34804 34432
rect 34820 34368 34884 34432
rect 34900 34368 34964 34432
rect 34980 34368 35044 34432
rect 35060 34368 35124 34432
rect 35140 34368 35204 34432
rect 35220 34368 35284 34432
rect 40740 34368 40804 34432
rect 40820 34368 40884 34432
rect 40900 34368 40964 34432
rect 40980 34368 41044 34432
rect 41060 34368 41124 34432
rect 41140 34368 41204 34432
rect 41220 34368 41284 34432
rect 46740 34368 46804 34432
rect 46820 34368 46884 34432
rect 46900 34368 46964 34432
rect 46980 34368 47044 34432
rect 47060 34368 47124 34432
rect 47140 34368 47204 34432
rect 47220 34368 47284 34432
rect 52740 34368 52804 34432
rect 52820 34368 52884 34432
rect 52900 34368 52964 34432
rect 52980 34368 53044 34432
rect 53060 34368 53124 34432
rect 53140 34368 53204 34432
rect 53220 34368 53284 34432
rect 58740 34368 58804 34432
rect 58820 34368 58884 34432
rect 58900 34368 58964 34432
rect 58980 34368 59044 34432
rect 59060 34368 59124 34432
rect 59140 34368 59204 34432
rect 59220 34368 59284 34432
rect 64740 34368 64804 34432
rect 64820 34368 64884 34432
rect 64900 34368 64964 34432
rect 64980 34368 65044 34432
rect 65060 34368 65124 34432
rect 65140 34368 65204 34432
rect 65220 34368 65284 34432
rect 70740 34368 70804 34432
rect 70820 34368 70884 34432
rect 70900 34368 70964 34432
rect 70980 34368 71044 34432
rect 71060 34368 71124 34432
rect 71140 34368 71204 34432
rect 71220 34368 71284 34432
rect 4740 34288 4804 34352
rect 4820 34288 4884 34352
rect 4900 34288 4964 34352
rect 4980 34288 5044 34352
rect 5060 34288 5124 34352
rect 5140 34288 5204 34352
rect 5220 34288 5284 34352
rect 10740 34288 10804 34352
rect 10820 34288 10884 34352
rect 10900 34288 10964 34352
rect 10980 34288 11044 34352
rect 11060 34288 11124 34352
rect 11140 34288 11204 34352
rect 11220 34288 11284 34352
rect 16740 34288 16804 34352
rect 16820 34288 16884 34352
rect 16900 34288 16964 34352
rect 16980 34288 17044 34352
rect 17060 34288 17124 34352
rect 17140 34288 17204 34352
rect 17220 34288 17284 34352
rect 22740 34288 22804 34352
rect 22820 34288 22884 34352
rect 22900 34288 22964 34352
rect 22980 34288 23044 34352
rect 23060 34288 23124 34352
rect 23140 34288 23204 34352
rect 23220 34288 23284 34352
rect 28740 34288 28804 34352
rect 28820 34288 28884 34352
rect 28900 34288 28964 34352
rect 28980 34288 29044 34352
rect 29060 34288 29124 34352
rect 29140 34288 29204 34352
rect 29220 34288 29284 34352
rect 34740 34288 34804 34352
rect 34820 34288 34884 34352
rect 34900 34288 34964 34352
rect 34980 34288 35044 34352
rect 35060 34288 35124 34352
rect 35140 34288 35204 34352
rect 35220 34288 35284 34352
rect 40740 34288 40804 34352
rect 40820 34288 40884 34352
rect 40900 34288 40964 34352
rect 40980 34288 41044 34352
rect 41060 34288 41124 34352
rect 41140 34288 41204 34352
rect 41220 34288 41284 34352
rect 46740 34288 46804 34352
rect 46820 34288 46884 34352
rect 46900 34288 46964 34352
rect 46980 34288 47044 34352
rect 47060 34288 47124 34352
rect 47140 34288 47204 34352
rect 47220 34288 47284 34352
rect 52740 34288 52804 34352
rect 52820 34288 52884 34352
rect 52900 34288 52964 34352
rect 52980 34288 53044 34352
rect 53060 34288 53124 34352
rect 53140 34288 53204 34352
rect 53220 34288 53284 34352
rect 58740 34288 58804 34352
rect 58820 34288 58884 34352
rect 58900 34288 58964 34352
rect 58980 34288 59044 34352
rect 59060 34288 59124 34352
rect 59140 34288 59204 34352
rect 59220 34288 59284 34352
rect 64740 34288 64804 34352
rect 64820 34288 64884 34352
rect 64900 34288 64964 34352
rect 64980 34288 65044 34352
rect 65060 34288 65124 34352
rect 65140 34288 65204 34352
rect 65220 34288 65284 34352
rect 70740 34288 70804 34352
rect 70820 34288 70884 34352
rect 70900 34288 70964 34352
rect 70980 34288 71044 34352
rect 71060 34288 71124 34352
rect 71140 34288 71204 34352
rect 71220 34288 71284 34352
rect 68508 33220 68572 33284
rect 1740 32176 1804 32240
rect 1820 32176 1884 32240
rect 1900 32176 1964 32240
rect 1980 32176 2044 32240
rect 2060 32176 2124 32240
rect 2140 32176 2204 32240
rect 2220 32176 2284 32240
rect 7740 32176 7804 32240
rect 7820 32176 7884 32240
rect 7900 32176 7964 32240
rect 7980 32176 8044 32240
rect 8060 32176 8124 32240
rect 8140 32176 8204 32240
rect 8220 32176 8284 32240
rect 13740 32176 13804 32240
rect 13820 32176 13884 32240
rect 13900 32176 13964 32240
rect 13980 32176 14044 32240
rect 14060 32176 14124 32240
rect 14140 32176 14204 32240
rect 14220 32176 14284 32240
rect 19740 32176 19804 32240
rect 19820 32176 19884 32240
rect 19900 32176 19964 32240
rect 19980 32176 20044 32240
rect 20060 32176 20124 32240
rect 20140 32176 20204 32240
rect 20220 32176 20284 32240
rect 25740 32176 25804 32240
rect 25820 32176 25884 32240
rect 25900 32176 25964 32240
rect 25980 32176 26044 32240
rect 26060 32176 26124 32240
rect 26140 32176 26204 32240
rect 26220 32176 26284 32240
rect 31740 32176 31804 32240
rect 31820 32176 31884 32240
rect 31900 32176 31964 32240
rect 31980 32176 32044 32240
rect 32060 32176 32124 32240
rect 32140 32176 32204 32240
rect 32220 32176 32284 32240
rect 37740 32176 37804 32240
rect 37820 32176 37884 32240
rect 37900 32176 37964 32240
rect 37980 32176 38044 32240
rect 38060 32176 38124 32240
rect 38140 32176 38204 32240
rect 38220 32176 38284 32240
rect 43740 32176 43804 32240
rect 43820 32176 43884 32240
rect 43900 32176 43964 32240
rect 43980 32176 44044 32240
rect 44060 32176 44124 32240
rect 44140 32176 44204 32240
rect 44220 32176 44284 32240
rect 49740 32176 49804 32240
rect 49820 32176 49884 32240
rect 49900 32176 49964 32240
rect 49980 32176 50044 32240
rect 50060 32176 50124 32240
rect 50140 32176 50204 32240
rect 50220 32176 50284 32240
rect 55740 32176 55804 32240
rect 55820 32176 55884 32240
rect 55900 32176 55964 32240
rect 55980 32176 56044 32240
rect 56060 32176 56124 32240
rect 56140 32176 56204 32240
rect 56220 32176 56284 32240
rect 61740 32176 61804 32240
rect 61820 32176 61884 32240
rect 61900 32176 61964 32240
rect 61980 32176 62044 32240
rect 62060 32176 62124 32240
rect 62140 32176 62204 32240
rect 62220 32176 62284 32240
rect 67740 32176 67804 32240
rect 67820 32176 67884 32240
rect 67900 32176 67964 32240
rect 67980 32176 68044 32240
rect 68060 32176 68124 32240
rect 68140 32176 68204 32240
rect 68220 32176 68284 32240
rect 73740 32176 73804 32240
rect 73820 32176 73884 32240
rect 73900 32176 73964 32240
rect 73980 32176 74044 32240
rect 74060 32176 74124 32240
rect 74140 32176 74204 32240
rect 74220 32176 74284 32240
rect 1740 32096 1804 32160
rect 1820 32096 1884 32160
rect 1900 32096 1964 32160
rect 1980 32096 2044 32160
rect 2060 32096 2124 32160
rect 2140 32096 2204 32160
rect 2220 32096 2284 32160
rect 7740 32096 7804 32160
rect 7820 32096 7884 32160
rect 7900 32096 7964 32160
rect 7980 32096 8044 32160
rect 8060 32096 8124 32160
rect 8140 32096 8204 32160
rect 8220 32096 8284 32160
rect 13740 32096 13804 32160
rect 13820 32096 13884 32160
rect 13900 32096 13964 32160
rect 13980 32096 14044 32160
rect 14060 32096 14124 32160
rect 14140 32096 14204 32160
rect 14220 32096 14284 32160
rect 19740 32096 19804 32160
rect 19820 32096 19884 32160
rect 19900 32096 19964 32160
rect 19980 32096 20044 32160
rect 20060 32096 20124 32160
rect 20140 32096 20204 32160
rect 20220 32096 20284 32160
rect 25740 32096 25804 32160
rect 25820 32096 25884 32160
rect 25900 32096 25964 32160
rect 25980 32096 26044 32160
rect 26060 32096 26124 32160
rect 26140 32096 26204 32160
rect 26220 32096 26284 32160
rect 31740 32096 31804 32160
rect 31820 32096 31884 32160
rect 31900 32096 31964 32160
rect 31980 32096 32044 32160
rect 32060 32096 32124 32160
rect 32140 32096 32204 32160
rect 32220 32096 32284 32160
rect 37740 32096 37804 32160
rect 37820 32096 37884 32160
rect 37900 32096 37964 32160
rect 37980 32096 38044 32160
rect 38060 32096 38124 32160
rect 38140 32096 38204 32160
rect 38220 32096 38284 32160
rect 43740 32096 43804 32160
rect 43820 32096 43884 32160
rect 43900 32096 43964 32160
rect 43980 32096 44044 32160
rect 44060 32096 44124 32160
rect 44140 32096 44204 32160
rect 44220 32096 44284 32160
rect 49740 32096 49804 32160
rect 49820 32096 49884 32160
rect 49900 32096 49964 32160
rect 49980 32096 50044 32160
rect 50060 32096 50124 32160
rect 50140 32096 50204 32160
rect 50220 32096 50284 32160
rect 55740 32096 55804 32160
rect 55820 32096 55884 32160
rect 55900 32096 55964 32160
rect 55980 32096 56044 32160
rect 56060 32096 56124 32160
rect 56140 32096 56204 32160
rect 56220 32096 56284 32160
rect 61740 32096 61804 32160
rect 61820 32096 61884 32160
rect 61900 32096 61964 32160
rect 61980 32096 62044 32160
rect 62060 32096 62124 32160
rect 62140 32096 62204 32160
rect 62220 32096 62284 32160
rect 67740 32096 67804 32160
rect 67820 32096 67884 32160
rect 67900 32096 67964 32160
rect 67980 32096 68044 32160
rect 68060 32096 68124 32160
rect 68140 32096 68204 32160
rect 68220 32096 68284 32160
rect 73740 32096 73804 32160
rect 73820 32096 73884 32160
rect 73900 32096 73964 32160
rect 73980 32096 74044 32160
rect 74060 32096 74124 32160
rect 74140 32096 74204 32160
rect 74220 32096 74284 32160
rect 1740 32016 1804 32080
rect 1820 32016 1884 32080
rect 1900 32016 1964 32080
rect 1980 32016 2044 32080
rect 2060 32016 2124 32080
rect 2140 32016 2204 32080
rect 2220 32016 2284 32080
rect 7740 32016 7804 32080
rect 7820 32016 7884 32080
rect 7900 32016 7964 32080
rect 7980 32016 8044 32080
rect 8060 32016 8124 32080
rect 8140 32016 8204 32080
rect 8220 32016 8284 32080
rect 13740 32016 13804 32080
rect 13820 32016 13884 32080
rect 13900 32016 13964 32080
rect 13980 32016 14044 32080
rect 14060 32016 14124 32080
rect 14140 32016 14204 32080
rect 14220 32016 14284 32080
rect 19740 32016 19804 32080
rect 19820 32016 19884 32080
rect 19900 32016 19964 32080
rect 19980 32016 20044 32080
rect 20060 32016 20124 32080
rect 20140 32016 20204 32080
rect 20220 32016 20284 32080
rect 25740 32016 25804 32080
rect 25820 32016 25884 32080
rect 25900 32016 25964 32080
rect 25980 32016 26044 32080
rect 26060 32016 26124 32080
rect 26140 32016 26204 32080
rect 26220 32016 26284 32080
rect 31740 32016 31804 32080
rect 31820 32016 31884 32080
rect 31900 32016 31964 32080
rect 31980 32016 32044 32080
rect 32060 32016 32124 32080
rect 32140 32016 32204 32080
rect 32220 32016 32284 32080
rect 37740 32016 37804 32080
rect 37820 32016 37884 32080
rect 37900 32016 37964 32080
rect 37980 32016 38044 32080
rect 38060 32016 38124 32080
rect 38140 32016 38204 32080
rect 38220 32016 38284 32080
rect 43740 32016 43804 32080
rect 43820 32016 43884 32080
rect 43900 32016 43964 32080
rect 43980 32016 44044 32080
rect 44060 32016 44124 32080
rect 44140 32016 44204 32080
rect 44220 32016 44284 32080
rect 49740 32016 49804 32080
rect 49820 32016 49884 32080
rect 49900 32016 49964 32080
rect 49980 32016 50044 32080
rect 50060 32016 50124 32080
rect 50140 32016 50204 32080
rect 50220 32016 50284 32080
rect 55740 32016 55804 32080
rect 55820 32016 55884 32080
rect 55900 32016 55964 32080
rect 55980 32016 56044 32080
rect 56060 32016 56124 32080
rect 56140 32016 56204 32080
rect 56220 32016 56284 32080
rect 61740 32016 61804 32080
rect 61820 32016 61884 32080
rect 61900 32016 61964 32080
rect 61980 32016 62044 32080
rect 62060 32016 62124 32080
rect 62140 32016 62204 32080
rect 62220 32016 62284 32080
rect 67740 32016 67804 32080
rect 67820 32016 67884 32080
rect 67900 32016 67964 32080
rect 67980 32016 68044 32080
rect 68060 32016 68124 32080
rect 68140 32016 68204 32080
rect 68220 32016 68284 32080
rect 73740 32016 73804 32080
rect 73820 32016 73884 32080
rect 73900 32016 73964 32080
rect 73980 32016 74044 32080
rect 74060 32016 74124 32080
rect 74140 32016 74204 32080
rect 74220 32016 74284 32080
rect 1740 31936 1804 32000
rect 1820 31936 1884 32000
rect 1900 31936 1964 32000
rect 1980 31936 2044 32000
rect 2060 31936 2124 32000
rect 2140 31936 2204 32000
rect 2220 31936 2284 32000
rect 7740 31936 7804 32000
rect 7820 31936 7884 32000
rect 7900 31936 7964 32000
rect 7980 31936 8044 32000
rect 8060 31936 8124 32000
rect 8140 31936 8204 32000
rect 8220 31936 8284 32000
rect 13740 31936 13804 32000
rect 13820 31936 13884 32000
rect 13900 31936 13964 32000
rect 13980 31936 14044 32000
rect 14060 31936 14124 32000
rect 14140 31936 14204 32000
rect 14220 31936 14284 32000
rect 19740 31936 19804 32000
rect 19820 31936 19884 32000
rect 19900 31936 19964 32000
rect 19980 31936 20044 32000
rect 20060 31936 20124 32000
rect 20140 31936 20204 32000
rect 20220 31936 20284 32000
rect 25740 31936 25804 32000
rect 25820 31936 25884 32000
rect 25900 31936 25964 32000
rect 25980 31936 26044 32000
rect 26060 31936 26124 32000
rect 26140 31936 26204 32000
rect 26220 31936 26284 32000
rect 31740 31936 31804 32000
rect 31820 31936 31884 32000
rect 31900 31936 31964 32000
rect 31980 31936 32044 32000
rect 32060 31936 32124 32000
rect 32140 31936 32204 32000
rect 32220 31936 32284 32000
rect 37740 31936 37804 32000
rect 37820 31936 37884 32000
rect 37900 31936 37964 32000
rect 37980 31936 38044 32000
rect 38060 31936 38124 32000
rect 38140 31936 38204 32000
rect 38220 31936 38284 32000
rect 43740 31936 43804 32000
rect 43820 31936 43884 32000
rect 43900 31936 43964 32000
rect 43980 31936 44044 32000
rect 44060 31936 44124 32000
rect 44140 31936 44204 32000
rect 44220 31936 44284 32000
rect 49740 31936 49804 32000
rect 49820 31936 49884 32000
rect 49900 31936 49964 32000
rect 49980 31936 50044 32000
rect 50060 31936 50124 32000
rect 50140 31936 50204 32000
rect 50220 31936 50284 32000
rect 55740 31936 55804 32000
rect 55820 31936 55884 32000
rect 55900 31936 55964 32000
rect 55980 31936 56044 32000
rect 56060 31936 56124 32000
rect 56140 31936 56204 32000
rect 56220 31936 56284 32000
rect 61740 31936 61804 32000
rect 61820 31936 61884 32000
rect 61900 31936 61964 32000
rect 61980 31936 62044 32000
rect 62060 31936 62124 32000
rect 62140 31936 62204 32000
rect 62220 31936 62284 32000
rect 67740 31936 67804 32000
rect 67820 31936 67884 32000
rect 67900 31936 67964 32000
rect 67980 31936 68044 32000
rect 68060 31936 68124 32000
rect 68140 31936 68204 32000
rect 68220 31936 68284 32000
rect 73740 31936 73804 32000
rect 73820 31936 73884 32000
rect 73900 31936 73964 32000
rect 73980 31936 74044 32000
rect 74060 31936 74124 32000
rect 74140 31936 74204 32000
rect 74220 31936 74284 32000
rect 67404 26480 67468 26484
rect 67404 26424 67418 26480
rect 67418 26424 67468 26480
rect 67404 26420 67468 26424
rect 63172 26148 63236 26212
rect 67404 26012 67468 26076
rect 4740 24528 4804 24592
rect 4820 24528 4884 24592
rect 4900 24528 4964 24592
rect 4980 24528 5044 24592
rect 5060 24528 5124 24592
rect 5140 24528 5204 24592
rect 5220 24528 5284 24592
rect 10740 24528 10804 24592
rect 10820 24528 10884 24592
rect 10900 24528 10964 24592
rect 10980 24528 11044 24592
rect 11060 24528 11124 24592
rect 11140 24528 11204 24592
rect 11220 24528 11284 24592
rect 16740 24528 16804 24592
rect 16820 24528 16884 24592
rect 16900 24528 16964 24592
rect 16980 24528 17044 24592
rect 17060 24528 17124 24592
rect 17140 24528 17204 24592
rect 17220 24528 17284 24592
rect 22740 24528 22804 24592
rect 22820 24528 22884 24592
rect 22900 24528 22964 24592
rect 22980 24528 23044 24592
rect 23060 24528 23124 24592
rect 23140 24528 23204 24592
rect 23220 24528 23284 24592
rect 28740 24528 28804 24592
rect 28820 24528 28884 24592
rect 28900 24528 28964 24592
rect 28980 24528 29044 24592
rect 29060 24528 29124 24592
rect 29140 24528 29204 24592
rect 29220 24528 29284 24592
rect 34740 24528 34804 24592
rect 34820 24528 34884 24592
rect 34900 24528 34964 24592
rect 34980 24528 35044 24592
rect 35060 24528 35124 24592
rect 35140 24528 35204 24592
rect 35220 24528 35284 24592
rect 40740 24528 40804 24592
rect 40820 24528 40884 24592
rect 40900 24528 40964 24592
rect 40980 24528 41044 24592
rect 41060 24528 41124 24592
rect 41140 24528 41204 24592
rect 41220 24528 41284 24592
rect 46740 24528 46804 24592
rect 46820 24528 46884 24592
rect 46900 24528 46964 24592
rect 46980 24528 47044 24592
rect 47060 24528 47124 24592
rect 47140 24528 47204 24592
rect 47220 24528 47284 24592
rect 52740 24528 52804 24592
rect 52820 24528 52884 24592
rect 52900 24528 52964 24592
rect 52980 24528 53044 24592
rect 53060 24528 53124 24592
rect 53140 24528 53204 24592
rect 53220 24528 53284 24592
rect 58740 24528 58804 24592
rect 58820 24528 58884 24592
rect 58900 24528 58964 24592
rect 58980 24528 59044 24592
rect 59060 24528 59124 24592
rect 59140 24528 59204 24592
rect 59220 24528 59284 24592
rect 64740 24528 64804 24592
rect 64820 24528 64884 24592
rect 64900 24528 64964 24592
rect 64980 24528 65044 24592
rect 65060 24528 65124 24592
rect 65140 24528 65204 24592
rect 65220 24528 65284 24592
rect 70740 24528 70804 24592
rect 70820 24528 70884 24592
rect 70900 24528 70964 24592
rect 70980 24528 71044 24592
rect 71060 24528 71124 24592
rect 71140 24528 71204 24592
rect 71220 24528 71284 24592
rect 4740 24448 4804 24512
rect 4820 24448 4884 24512
rect 4900 24448 4964 24512
rect 4980 24448 5044 24512
rect 5060 24448 5124 24512
rect 5140 24448 5204 24512
rect 5220 24448 5284 24512
rect 10740 24448 10804 24512
rect 10820 24448 10884 24512
rect 10900 24448 10964 24512
rect 10980 24448 11044 24512
rect 11060 24448 11124 24512
rect 11140 24448 11204 24512
rect 11220 24448 11284 24512
rect 16740 24448 16804 24512
rect 16820 24448 16884 24512
rect 16900 24448 16964 24512
rect 16980 24448 17044 24512
rect 17060 24448 17124 24512
rect 17140 24448 17204 24512
rect 17220 24448 17284 24512
rect 22740 24448 22804 24512
rect 22820 24448 22884 24512
rect 22900 24448 22964 24512
rect 22980 24448 23044 24512
rect 23060 24448 23124 24512
rect 23140 24448 23204 24512
rect 23220 24448 23284 24512
rect 28740 24448 28804 24512
rect 28820 24448 28884 24512
rect 28900 24448 28964 24512
rect 28980 24448 29044 24512
rect 29060 24448 29124 24512
rect 29140 24448 29204 24512
rect 29220 24448 29284 24512
rect 34740 24448 34804 24512
rect 34820 24448 34884 24512
rect 34900 24448 34964 24512
rect 34980 24448 35044 24512
rect 35060 24448 35124 24512
rect 35140 24448 35204 24512
rect 35220 24448 35284 24512
rect 40740 24448 40804 24512
rect 40820 24448 40884 24512
rect 40900 24448 40964 24512
rect 40980 24448 41044 24512
rect 41060 24448 41124 24512
rect 41140 24448 41204 24512
rect 41220 24448 41284 24512
rect 46740 24448 46804 24512
rect 46820 24448 46884 24512
rect 46900 24448 46964 24512
rect 46980 24448 47044 24512
rect 47060 24448 47124 24512
rect 47140 24448 47204 24512
rect 47220 24448 47284 24512
rect 52740 24448 52804 24512
rect 52820 24448 52884 24512
rect 52900 24448 52964 24512
rect 52980 24448 53044 24512
rect 53060 24448 53124 24512
rect 53140 24448 53204 24512
rect 53220 24448 53284 24512
rect 58740 24448 58804 24512
rect 58820 24448 58884 24512
rect 58900 24448 58964 24512
rect 58980 24448 59044 24512
rect 59060 24448 59124 24512
rect 59140 24448 59204 24512
rect 59220 24448 59284 24512
rect 64740 24448 64804 24512
rect 64820 24448 64884 24512
rect 64900 24448 64964 24512
rect 64980 24448 65044 24512
rect 65060 24448 65124 24512
rect 65140 24448 65204 24512
rect 65220 24448 65284 24512
rect 70740 24448 70804 24512
rect 70820 24448 70884 24512
rect 70900 24448 70964 24512
rect 70980 24448 71044 24512
rect 71060 24448 71124 24512
rect 71140 24448 71204 24512
rect 71220 24448 71284 24512
rect 4740 24368 4804 24432
rect 4820 24368 4884 24432
rect 4900 24368 4964 24432
rect 4980 24368 5044 24432
rect 5060 24368 5124 24432
rect 5140 24368 5204 24432
rect 5220 24368 5284 24432
rect 10740 24368 10804 24432
rect 10820 24368 10884 24432
rect 10900 24368 10964 24432
rect 10980 24368 11044 24432
rect 11060 24368 11124 24432
rect 11140 24368 11204 24432
rect 11220 24368 11284 24432
rect 16740 24368 16804 24432
rect 16820 24368 16884 24432
rect 16900 24368 16964 24432
rect 16980 24368 17044 24432
rect 17060 24368 17124 24432
rect 17140 24368 17204 24432
rect 17220 24368 17284 24432
rect 22740 24368 22804 24432
rect 22820 24368 22884 24432
rect 22900 24368 22964 24432
rect 22980 24368 23044 24432
rect 23060 24368 23124 24432
rect 23140 24368 23204 24432
rect 23220 24368 23284 24432
rect 28740 24368 28804 24432
rect 28820 24368 28884 24432
rect 28900 24368 28964 24432
rect 28980 24368 29044 24432
rect 29060 24368 29124 24432
rect 29140 24368 29204 24432
rect 29220 24368 29284 24432
rect 34740 24368 34804 24432
rect 34820 24368 34884 24432
rect 34900 24368 34964 24432
rect 34980 24368 35044 24432
rect 35060 24368 35124 24432
rect 35140 24368 35204 24432
rect 35220 24368 35284 24432
rect 40740 24368 40804 24432
rect 40820 24368 40884 24432
rect 40900 24368 40964 24432
rect 40980 24368 41044 24432
rect 41060 24368 41124 24432
rect 41140 24368 41204 24432
rect 41220 24368 41284 24432
rect 46740 24368 46804 24432
rect 46820 24368 46884 24432
rect 46900 24368 46964 24432
rect 46980 24368 47044 24432
rect 47060 24368 47124 24432
rect 47140 24368 47204 24432
rect 47220 24368 47284 24432
rect 52740 24368 52804 24432
rect 52820 24368 52884 24432
rect 52900 24368 52964 24432
rect 52980 24368 53044 24432
rect 53060 24368 53124 24432
rect 53140 24368 53204 24432
rect 53220 24368 53284 24432
rect 58740 24368 58804 24432
rect 58820 24368 58884 24432
rect 58900 24368 58964 24432
rect 58980 24368 59044 24432
rect 59060 24368 59124 24432
rect 59140 24368 59204 24432
rect 59220 24368 59284 24432
rect 64740 24368 64804 24432
rect 64820 24368 64884 24432
rect 64900 24368 64964 24432
rect 64980 24368 65044 24432
rect 65060 24368 65124 24432
rect 65140 24368 65204 24432
rect 65220 24368 65284 24432
rect 70740 24368 70804 24432
rect 70820 24368 70884 24432
rect 70900 24368 70964 24432
rect 70980 24368 71044 24432
rect 71060 24368 71124 24432
rect 71140 24368 71204 24432
rect 71220 24368 71284 24432
rect 4740 24288 4804 24352
rect 4820 24288 4884 24352
rect 4900 24288 4964 24352
rect 4980 24288 5044 24352
rect 5060 24288 5124 24352
rect 5140 24288 5204 24352
rect 5220 24288 5284 24352
rect 10740 24288 10804 24352
rect 10820 24288 10884 24352
rect 10900 24288 10964 24352
rect 10980 24288 11044 24352
rect 11060 24288 11124 24352
rect 11140 24288 11204 24352
rect 11220 24288 11284 24352
rect 16740 24288 16804 24352
rect 16820 24288 16884 24352
rect 16900 24288 16964 24352
rect 16980 24288 17044 24352
rect 17060 24288 17124 24352
rect 17140 24288 17204 24352
rect 17220 24288 17284 24352
rect 22740 24288 22804 24352
rect 22820 24288 22884 24352
rect 22900 24288 22964 24352
rect 22980 24288 23044 24352
rect 23060 24288 23124 24352
rect 23140 24288 23204 24352
rect 23220 24288 23284 24352
rect 28740 24288 28804 24352
rect 28820 24288 28884 24352
rect 28900 24288 28964 24352
rect 28980 24288 29044 24352
rect 29060 24288 29124 24352
rect 29140 24288 29204 24352
rect 29220 24288 29284 24352
rect 34740 24288 34804 24352
rect 34820 24288 34884 24352
rect 34900 24288 34964 24352
rect 34980 24288 35044 24352
rect 35060 24288 35124 24352
rect 35140 24288 35204 24352
rect 35220 24288 35284 24352
rect 40740 24288 40804 24352
rect 40820 24288 40884 24352
rect 40900 24288 40964 24352
rect 40980 24288 41044 24352
rect 41060 24288 41124 24352
rect 41140 24288 41204 24352
rect 41220 24288 41284 24352
rect 46740 24288 46804 24352
rect 46820 24288 46884 24352
rect 46900 24288 46964 24352
rect 46980 24288 47044 24352
rect 47060 24288 47124 24352
rect 47140 24288 47204 24352
rect 47220 24288 47284 24352
rect 52740 24288 52804 24352
rect 52820 24288 52884 24352
rect 52900 24288 52964 24352
rect 52980 24288 53044 24352
rect 53060 24288 53124 24352
rect 53140 24288 53204 24352
rect 53220 24288 53284 24352
rect 58740 24288 58804 24352
rect 58820 24288 58884 24352
rect 58900 24288 58964 24352
rect 58980 24288 59044 24352
rect 59060 24288 59124 24352
rect 59140 24288 59204 24352
rect 59220 24288 59284 24352
rect 64740 24288 64804 24352
rect 64820 24288 64884 24352
rect 64900 24288 64964 24352
rect 64980 24288 65044 24352
rect 65060 24288 65124 24352
rect 65140 24288 65204 24352
rect 65220 24288 65284 24352
rect 70740 24288 70804 24352
rect 70820 24288 70884 24352
rect 70900 24288 70964 24352
rect 70980 24288 71044 24352
rect 71060 24288 71124 24352
rect 71140 24288 71204 24352
rect 71220 24288 71284 24352
rect 66484 23564 66548 23628
rect 66300 23428 66364 23492
rect 66668 22340 66732 22404
rect 1740 22176 1804 22240
rect 1820 22176 1884 22240
rect 1900 22176 1964 22240
rect 1980 22176 2044 22240
rect 2060 22176 2124 22240
rect 2140 22176 2204 22240
rect 2220 22176 2284 22240
rect 7740 22176 7804 22240
rect 7820 22176 7884 22240
rect 7900 22176 7964 22240
rect 7980 22176 8044 22240
rect 8060 22176 8124 22240
rect 8140 22176 8204 22240
rect 8220 22176 8284 22240
rect 13740 22176 13804 22240
rect 13820 22176 13884 22240
rect 13900 22176 13964 22240
rect 13980 22176 14044 22240
rect 14060 22176 14124 22240
rect 14140 22176 14204 22240
rect 14220 22176 14284 22240
rect 19740 22176 19804 22240
rect 19820 22176 19884 22240
rect 19900 22176 19964 22240
rect 19980 22176 20044 22240
rect 20060 22176 20124 22240
rect 20140 22176 20204 22240
rect 20220 22176 20284 22240
rect 25740 22176 25804 22240
rect 25820 22176 25884 22240
rect 25900 22176 25964 22240
rect 25980 22176 26044 22240
rect 26060 22176 26124 22240
rect 26140 22176 26204 22240
rect 26220 22176 26284 22240
rect 31740 22176 31804 22240
rect 31820 22176 31884 22240
rect 31900 22176 31964 22240
rect 31980 22176 32044 22240
rect 32060 22176 32124 22240
rect 32140 22176 32204 22240
rect 32220 22176 32284 22240
rect 37740 22176 37804 22240
rect 37820 22176 37884 22240
rect 37900 22176 37964 22240
rect 37980 22176 38044 22240
rect 38060 22176 38124 22240
rect 38140 22176 38204 22240
rect 38220 22176 38284 22240
rect 43740 22176 43804 22240
rect 43820 22176 43884 22240
rect 43900 22176 43964 22240
rect 43980 22176 44044 22240
rect 44060 22176 44124 22240
rect 44140 22176 44204 22240
rect 44220 22176 44284 22240
rect 49740 22176 49804 22240
rect 49820 22176 49884 22240
rect 49900 22176 49964 22240
rect 49980 22176 50044 22240
rect 50060 22176 50124 22240
rect 50140 22176 50204 22240
rect 50220 22176 50284 22240
rect 55740 22176 55804 22240
rect 55820 22176 55884 22240
rect 55900 22176 55964 22240
rect 55980 22176 56044 22240
rect 56060 22176 56124 22240
rect 56140 22176 56204 22240
rect 56220 22176 56284 22240
rect 61740 22176 61804 22240
rect 61820 22176 61884 22240
rect 61900 22176 61964 22240
rect 61980 22176 62044 22240
rect 62060 22176 62124 22240
rect 62140 22176 62204 22240
rect 62220 22176 62284 22240
rect 67740 22176 67804 22240
rect 67820 22176 67884 22240
rect 67900 22176 67964 22240
rect 67980 22176 68044 22240
rect 68060 22176 68124 22240
rect 68140 22176 68204 22240
rect 68220 22176 68284 22240
rect 73740 22176 73804 22240
rect 73820 22176 73884 22240
rect 73900 22176 73964 22240
rect 73980 22176 74044 22240
rect 74060 22176 74124 22240
rect 74140 22176 74204 22240
rect 74220 22176 74284 22240
rect 1740 22096 1804 22160
rect 1820 22096 1884 22160
rect 1900 22096 1964 22160
rect 1980 22096 2044 22160
rect 2060 22096 2124 22160
rect 2140 22096 2204 22160
rect 2220 22096 2284 22160
rect 7740 22096 7804 22160
rect 7820 22096 7884 22160
rect 7900 22096 7964 22160
rect 7980 22096 8044 22160
rect 8060 22096 8124 22160
rect 8140 22096 8204 22160
rect 8220 22096 8284 22160
rect 13740 22096 13804 22160
rect 13820 22096 13884 22160
rect 13900 22096 13964 22160
rect 13980 22096 14044 22160
rect 14060 22096 14124 22160
rect 14140 22096 14204 22160
rect 14220 22096 14284 22160
rect 19740 22096 19804 22160
rect 19820 22096 19884 22160
rect 19900 22096 19964 22160
rect 19980 22096 20044 22160
rect 20060 22096 20124 22160
rect 20140 22096 20204 22160
rect 20220 22096 20284 22160
rect 25740 22096 25804 22160
rect 25820 22096 25884 22160
rect 25900 22096 25964 22160
rect 25980 22096 26044 22160
rect 26060 22096 26124 22160
rect 26140 22096 26204 22160
rect 26220 22096 26284 22160
rect 31740 22096 31804 22160
rect 31820 22096 31884 22160
rect 31900 22096 31964 22160
rect 31980 22096 32044 22160
rect 32060 22096 32124 22160
rect 32140 22096 32204 22160
rect 32220 22096 32284 22160
rect 37740 22096 37804 22160
rect 37820 22096 37884 22160
rect 37900 22096 37964 22160
rect 37980 22096 38044 22160
rect 38060 22096 38124 22160
rect 38140 22096 38204 22160
rect 38220 22096 38284 22160
rect 43740 22096 43804 22160
rect 43820 22096 43884 22160
rect 43900 22096 43964 22160
rect 43980 22096 44044 22160
rect 44060 22096 44124 22160
rect 44140 22096 44204 22160
rect 44220 22096 44284 22160
rect 49740 22096 49804 22160
rect 49820 22096 49884 22160
rect 49900 22096 49964 22160
rect 49980 22096 50044 22160
rect 50060 22096 50124 22160
rect 50140 22096 50204 22160
rect 50220 22096 50284 22160
rect 55740 22096 55804 22160
rect 55820 22096 55884 22160
rect 55900 22096 55964 22160
rect 55980 22096 56044 22160
rect 56060 22096 56124 22160
rect 56140 22096 56204 22160
rect 56220 22096 56284 22160
rect 61740 22096 61804 22160
rect 61820 22096 61884 22160
rect 61900 22096 61964 22160
rect 61980 22096 62044 22160
rect 62060 22096 62124 22160
rect 62140 22096 62204 22160
rect 62220 22096 62284 22160
rect 67740 22096 67804 22160
rect 67820 22096 67884 22160
rect 67900 22096 67964 22160
rect 67980 22096 68044 22160
rect 68060 22096 68124 22160
rect 68140 22096 68204 22160
rect 68220 22096 68284 22160
rect 73740 22096 73804 22160
rect 73820 22096 73884 22160
rect 73900 22096 73964 22160
rect 73980 22096 74044 22160
rect 74060 22096 74124 22160
rect 74140 22096 74204 22160
rect 74220 22096 74284 22160
rect 1740 22016 1804 22080
rect 1820 22016 1884 22080
rect 1900 22016 1964 22080
rect 1980 22016 2044 22080
rect 2060 22016 2124 22080
rect 2140 22016 2204 22080
rect 2220 22016 2284 22080
rect 7740 22016 7804 22080
rect 7820 22016 7884 22080
rect 7900 22016 7964 22080
rect 7980 22016 8044 22080
rect 8060 22016 8124 22080
rect 8140 22016 8204 22080
rect 8220 22016 8284 22080
rect 13740 22016 13804 22080
rect 13820 22016 13884 22080
rect 13900 22016 13964 22080
rect 13980 22016 14044 22080
rect 14060 22016 14124 22080
rect 14140 22016 14204 22080
rect 14220 22016 14284 22080
rect 19740 22016 19804 22080
rect 19820 22016 19884 22080
rect 19900 22016 19964 22080
rect 19980 22016 20044 22080
rect 20060 22016 20124 22080
rect 20140 22016 20204 22080
rect 20220 22016 20284 22080
rect 25740 22016 25804 22080
rect 25820 22016 25884 22080
rect 25900 22016 25964 22080
rect 25980 22016 26044 22080
rect 26060 22016 26124 22080
rect 26140 22016 26204 22080
rect 26220 22016 26284 22080
rect 31740 22016 31804 22080
rect 31820 22016 31884 22080
rect 31900 22016 31964 22080
rect 31980 22016 32044 22080
rect 32060 22016 32124 22080
rect 32140 22016 32204 22080
rect 32220 22016 32284 22080
rect 37740 22016 37804 22080
rect 37820 22016 37884 22080
rect 37900 22016 37964 22080
rect 37980 22016 38044 22080
rect 38060 22016 38124 22080
rect 38140 22016 38204 22080
rect 38220 22016 38284 22080
rect 43740 22016 43804 22080
rect 43820 22016 43884 22080
rect 43900 22016 43964 22080
rect 43980 22016 44044 22080
rect 44060 22016 44124 22080
rect 44140 22016 44204 22080
rect 44220 22016 44284 22080
rect 49740 22016 49804 22080
rect 49820 22016 49884 22080
rect 49900 22016 49964 22080
rect 49980 22016 50044 22080
rect 50060 22016 50124 22080
rect 50140 22016 50204 22080
rect 50220 22016 50284 22080
rect 55740 22016 55804 22080
rect 55820 22016 55884 22080
rect 55900 22016 55964 22080
rect 55980 22016 56044 22080
rect 56060 22016 56124 22080
rect 56140 22016 56204 22080
rect 56220 22016 56284 22080
rect 61740 22016 61804 22080
rect 61820 22016 61884 22080
rect 61900 22016 61964 22080
rect 61980 22016 62044 22080
rect 62060 22016 62124 22080
rect 62140 22016 62204 22080
rect 62220 22016 62284 22080
rect 67740 22016 67804 22080
rect 67820 22016 67884 22080
rect 67900 22016 67964 22080
rect 67980 22016 68044 22080
rect 68060 22016 68124 22080
rect 68140 22016 68204 22080
rect 68220 22016 68284 22080
rect 73740 22016 73804 22080
rect 73820 22016 73884 22080
rect 73900 22016 73964 22080
rect 73980 22016 74044 22080
rect 74060 22016 74124 22080
rect 74140 22016 74204 22080
rect 74220 22016 74284 22080
rect 1740 21936 1804 22000
rect 1820 21936 1884 22000
rect 1900 21936 1964 22000
rect 1980 21936 2044 22000
rect 2060 21936 2124 22000
rect 2140 21936 2204 22000
rect 2220 21936 2284 22000
rect 7740 21936 7804 22000
rect 7820 21936 7884 22000
rect 7900 21936 7964 22000
rect 7980 21936 8044 22000
rect 8060 21936 8124 22000
rect 8140 21936 8204 22000
rect 8220 21936 8284 22000
rect 13740 21936 13804 22000
rect 13820 21936 13884 22000
rect 13900 21936 13964 22000
rect 13980 21936 14044 22000
rect 14060 21936 14124 22000
rect 14140 21936 14204 22000
rect 14220 21936 14284 22000
rect 19740 21936 19804 22000
rect 19820 21936 19884 22000
rect 19900 21936 19964 22000
rect 19980 21936 20044 22000
rect 20060 21936 20124 22000
rect 20140 21936 20204 22000
rect 20220 21936 20284 22000
rect 25740 21936 25804 22000
rect 25820 21936 25884 22000
rect 25900 21936 25964 22000
rect 25980 21936 26044 22000
rect 26060 21936 26124 22000
rect 26140 21936 26204 22000
rect 26220 21936 26284 22000
rect 31740 21936 31804 22000
rect 31820 21936 31884 22000
rect 31900 21936 31964 22000
rect 31980 21936 32044 22000
rect 32060 21936 32124 22000
rect 32140 21936 32204 22000
rect 32220 21936 32284 22000
rect 37740 21936 37804 22000
rect 37820 21936 37884 22000
rect 37900 21936 37964 22000
rect 37980 21936 38044 22000
rect 38060 21936 38124 22000
rect 38140 21936 38204 22000
rect 38220 21936 38284 22000
rect 43740 21936 43804 22000
rect 43820 21936 43884 22000
rect 43900 21936 43964 22000
rect 43980 21936 44044 22000
rect 44060 21936 44124 22000
rect 44140 21936 44204 22000
rect 44220 21936 44284 22000
rect 49740 21936 49804 22000
rect 49820 21936 49884 22000
rect 49900 21936 49964 22000
rect 49980 21936 50044 22000
rect 50060 21936 50124 22000
rect 50140 21936 50204 22000
rect 50220 21936 50284 22000
rect 55740 21936 55804 22000
rect 55820 21936 55884 22000
rect 55900 21936 55964 22000
rect 55980 21936 56044 22000
rect 56060 21936 56124 22000
rect 56140 21936 56204 22000
rect 56220 21936 56284 22000
rect 61740 21936 61804 22000
rect 61820 21936 61884 22000
rect 61900 21936 61964 22000
rect 61980 21936 62044 22000
rect 62060 21936 62124 22000
rect 62140 21936 62204 22000
rect 62220 21936 62284 22000
rect 67740 21936 67804 22000
rect 67820 21936 67884 22000
rect 67900 21936 67964 22000
rect 67980 21936 68044 22000
rect 68060 21936 68124 22000
rect 68140 21936 68204 22000
rect 68220 21936 68284 22000
rect 73740 21936 73804 22000
rect 73820 21936 73884 22000
rect 73900 21936 73964 22000
rect 73980 21936 74044 22000
rect 74060 21936 74124 22000
rect 74140 21936 74204 22000
rect 74220 21936 74284 22000
rect 63540 16492 63604 16556
rect 63724 14724 63788 14788
rect 64460 14724 64524 14788
rect 4740 14528 4804 14592
rect 4820 14528 4884 14592
rect 4900 14528 4964 14592
rect 4980 14528 5044 14592
rect 5060 14528 5124 14592
rect 5140 14528 5204 14592
rect 5220 14528 5284 14592
rect 10740 14528 10804 14592
rect 10820 14528 10884 14592
rect 10900 14528 10964 14592
rect 10980 14528 11044 14592
rect 11060 14528 11124 14592
rect 11140 14528 11204 14592
rect 11220 14528 11284 14592
rect 16740 14528 16804 14592
rect 16820 14528 16884 14592
rect 16900 14528 16964 14592
rect 16980 14528 17044 14592
rect 17060 14528 17124 14592
rect 17140 14528 17204 14592
rect 17220 14528 17284 14592
rect 22740 14528 22804 14592
rect 22820 14528 22884 14592
rect 22900 14528 22964 14592
rect 22980 14528 23044 14592
rect 23060 14528 23124 14592
rect 23140 14528 23204 14592
rect 23220 14528 23284 14592
rect 28740 14528 28804 14592
rect 28820 14528 28884 14592
rect 28900 14528 28964 14592
rect 28980 14528 29044 14592
rect 29060 14528 29124 14592
rect 29140 14528 29204 14592
rect 29220 14528 29284 14592
rect 34740 14528 34804 14592
rect 34820 14528 34884 14592
rect 34900 14528 34964 14592
rect 34980 14528 35044 14592
rect 35060 14528 35124 14592
rect 35140 14528 35204 14592
rect 35220 14528 35284 14592
rect 40740 14528 40804 14592
rect 40820 14528 40884 14592
rect 40900 14528 40964 14592
rect 40980 14528 41044 14592
rect 41060 14528 41124 14592
rect 41140 14528 41204 14592
rect 41220 14528 41284 14592
rect 46740 14528 46804 14592
rect 46820 14528 46884 14592
rect 46900 14528 46964 14592
rect 46980 14528 47044 14592
rect 47060 14528 47124 14592
rect 47140 14528 47204 14592
rect 47220 14528 47284 14592
rect 52740 14528 52804 14592
rect 52820 14528 52884 14592
rect 52900 14528 52964 14592
rect 52980 14528 53044 14592
rect 53060 14528 53124 14592
rect 53140 14528 53204 14592
rect 53220 14528 53284 14592
rect 58740 14528 58804 14592
rect 58820 14528 58884 14592
rect 58900 14528 58964 14592
rect 58980 14528 59044 14592
rect 59060 14528 59124 14592
rect 59140 14528 59204 14592
rect 59220 14528 59284 14592
rect 64740 14528 64804 14592
rect 64820 14528 64884 14592
rect 64900 14528 64964 14592
rect 64980 14528 65044 14592
rect 65060 14528 65124 14592
rect 65140 14528 65204 14592
rect 65220 14528 65284 14592
rect 70740 14528 70804 14592
rect 70820 14528 70884 14592
rect 70900 14528 70964 14592
rect 70980 14528 71044 14592
rect 71060 14528 71124 14592
rect 71140 14528 71204 14592
rect 71220 14528 71284 14592
rect 4740 14448 4804 14512
rect 4820 14448 4884 14512
rect 4900 14448 4964 14512
rect 4980 14448 5044 14512
rect 5060 14448 5124 14512
rect 5140 14448 5204 14512
rect 5220 14448 5284 14512
rect 10740 14448 10804 14512
rect 10820 14448 10884 14512
rect 10900 14448 10964 14512
rect 10980 14448 11044 14512
rect 11060 14448 11124 14512
rect 11140 14448 11204 14512
rect 11220 14448 11284 14512
rect 16740 14448 16804 14512
rect 16820 14448 16884 14512
rect 16900 14448 16964 14512
rect 16980 14448 17044 14512
rect 17060 14448 17124 14512
rect 17140 14448 17204 14512
rect 17220 14448 17284 14512
rect 22740 14448 22804 14512
rect 22820 14448 22884 14512
rect 22900 14448 22964 14512
rect 22980 14448 23044 14512
rect 23060 14448 23124 14512
rect 23140 14448 23204 14512
rect 23220 14448 23284 14512
rect 28740 14448 28804 14512
rect 28820 14448 28884 14512
rect 28900 14448 28964 14512
rect 28980 14448 29044 14512
rect 29060 14448 29124 14512
rect 29140 14448 29204 14512
rect 29220 14448 29284 14512
rect 34740 14448 34804 14512
rect 34820 14448 34884 14512
rect 34900 14448 34964 14512
rect 34980 14448 35044 14512
rect 35060 14448 35124 14512
rect 35140 14448 35204 14512
rect 35220 14448 35284 14512
rect 40740 14448 40804 14512
rect 40820 14448 40884 14512
rect 40900 14448 40964 14512
rect 40980 14448 41044 14512
rect 41060 14448 41124 14512
rect 41140 14448 41204 14512
rect 41220 14448 41284 14512
rect 46740 14448 46804 14512
rect 46820 14448 46884 14512
rect 46900 14448 46964 14512
rect 46980 14448 47044 14512
rect 47060 14448 47124 14512
rect 47140 14448 47204 14512
rect 47220 14448 47284 14512
rect 52740 14448 52804 14512
rect 52820 14448 52884 14512
rect 52900 14448 52964 14512
rect 52980 14448 53044 14512
rect 53060 14448 53124 14512
rect 53140 14448 53204 14512
rect 53220 14448 53284 14512
rect 58740 14448 58804 14512
rect 58820 14448 58884 14512
rect 58900 14448 58964 14512
rect 58980 14448 59044 14512
rect 59060 14448 59124 14512
rect 59140 14448 59204 14512
rect 59220 14448 59284 14512
rect 64740 14448 64804 14512
rect 64820 14448 64884 14512
rect 64900 14448 64964 14512
rect 64980 14448 65044 14512
rect 65060 14448 65124 14512
rect 65140 14448 65204 14512
rect 65220 14448 65284 14512
rect 70740 14448 70804 14512
rect 70820 14448 70884 14512
rect 70900 14448 70964 14512
rect 70980 14448 71044 14512
rect 71060 14448 71124 14512
rect 71140 14448 71204 14512
rect 71220 14448 71284 14512
rect 4740 14368 4804 14432
rect 4820 14368 4884 14432
rect 4900 14368 4964 14432
rect 4980 14368 5044 14432
rect 5060 14368 5124 14432
rect 5140 14368 5204 14432
rect 5220 14368 5284 14432
rect 10740 14368 10804 14432
rect 10820 14368 10884 14432
rect 10900 14368 10964 14432
rect 10980 14368 11044 14432
rect 11060 14368 11124 14432
rect 11140 14368 11204 14432
rect 11220 14368 11284 14432
rect 16740 14368 16804 14432
rect 16820 14368 16884 14432
rect 16900 14368 16964 14432
rect 16980 14368 17044 14432
rect 17060 14368 17124 14432
rect 17140 14368 17204 14432
rect 17220 14368 17284 14432
rect 22740 14368 22804 14432
rect 22820 14368 22884 14432
rect 22900 14368 22964 14432
rect 22980 14368 23044 14432
rect 23060 14368 23124 14432
rect 23140 14368 23204 14432
rect 23220 14368 23284 14432
rect 28740 14368 28804 14432
rect 28820 14368 28884 14432
rect 28900 14368 28964 14432
rect 28980 14368 29044 14432
rect 29060 14368 29124 14432
rect 29140 14368 29204 14432
rect 29220 14368 29284 14432
rect 34740 14368 34804 14432
rect 34820 14368 34884 14432
rect 34900 14368 34964 14432
rect 34980 14368 35044 14432
rect 35060 14368 35124 14432
rect 35140 14368 35204 14432
rect 35220 14368 35284 14432
rect 40740 14368 40804 14432
rect 40820 14368 40884 14432
rect 40900 14368 40964 14432
rect 40980 14368 41044 14432
rect 41060 14368 41124 14432
rect 41140 14368 41204 14432
rect 41220 14368 41284 14432
rect 46740 14368 46804 14432
rect 46820 14368 46884 14432
rect 46900 14368 46964 14432
rect 46980 14368 47044 14432
rect 47060 14368 47124 14432
rect 47140 14368 47204 14432
rect 47220 14368 47284 14432
rect 52740 14368 52804 14432
rect 52820 14368 52884 14432
rect 52900 14368 52964 14432
rect 52980 14368 53044 14432
rect 53060 14368 53124 14432
rect 53140 14368 53204 14432
rect 53220 14368 53284 14432
rect 58740 14368 58804 14432
rect 58820 14368 58884 14432
rect 58900 14368 58964 14432
rect 58980 14368 59044 14432
rect 59060 14368 59124 14432
rect 59140 14368 59204 14432
rect 59220 14368 59284 14432
rect 64740 14368 64804 14432
rect 64820 14368 64884 14432
rect 64900 14368 64964 14432
rect 64980 14368 65044 14432
rect 65060 14368 65124 14432
rect 65140 14368 65204 14432
rect 65220 14368 65284 14432
rect 70740 14368 70804 14432
rect 70820 14368 70884 14432
rect 70900 14368 70964 14432
rect 70980 14368 71044 14432
rect 71060 14368 71124 14432
rect 71140 14368 71204 14432
rect 71220 14368 71284 14432
rect 4740 14288 4804 14352
rect 4820 14288 4884 14352
rect 4900 14288 4964 14352
rect 4980 14288 5044 14352
rect 5060 14288 5124 14352
rect 5140 14288 5204 14352
rect 5220 14288 5284 14352
rect 10740 14288 10804 14352
rect 10820 14288 10884 14352
rect 10900 14288 10964 14352
rect 10980 14288 11044 14352
rect 11060 14288 11124 14352
rect 11140 14288 11204 14352
rect 11220 14288 11284 14352
rect 16740 14288 16804 14352
rect 16820 14288 16884 14352
rect 16900 14288 16964 14352
rect 16980 14288 17044 14352
rect 17060 14288 17124 14352
rect 17140 14288 17204 14352
rect 17220 14288 17284 14352
rect 22740 14288 22804 14352
rect 22820 14288 22884 14352
rect 22900 14288 22964 14352
rect 22980 14288 23044 14352
rect 23060 14288 23124 14352
rect 23140 14288 23204 14352
rect 23220 14288 23284 14352
rect 28740 14288 28804 14352
rect 28820 14288 28884 14352
rect 28900 14288 28964 14352
rect 28980 14288 29044 14352
rect 29060 14288 29124 14352
rect 29140 14288 29204 14352
rect 29220 14288 29284 14352
rect 34740 14288 34804 14352
rect 34820 14288 34884 14352
rect 34900 14288 34964 14352
rect 34980 14288 35044 14352
rect 35060 14288 35124 14352
rect 35140 14288 35204 14352
rect 35220 14288 35284 14352
rect 40740 14288 40804 14352
rect 40820 14288 40884 14352
rect 40900 14288 40964 14352
rect 40980 14288 41044 14352
rect 41060 14288 41124 14352
rect 41140 14288 41204 14352
rect 41220 14288 41284 14352
rect 46740 14288 46804 14352
rect 46820 14288 46884 14352
rect 46900 14288 46964 14352
rect 46980 14288 47044 14352
rect 47060 14288 47124 14352
rect 47140 14288 47204 14352
rect 47220 14288 47284 14352
rect 52740 14288 52804 14352
rect 52820 14288 52884 14352
rect 52900 14288 52964 14352
rect 52980 14288 53044 14352
rect 53060 14288 53124 14352
rect 53140 14288 53204 14352
rect 53220 14288 53284 14352
rect 58740 14288 58804 14352
rect 58820 14288 58884 14352
rect 58900 14288 58964 14352
rect 58980 14288 59044 14352
rect 59060 14288 59124 14352
rect 59140 14288 59204 14352
rect 59220 14288 59284 14352
rect 64740 14288 64804 14352
rect 64820 14288 64884 14352
rect 64900 14288 64964 14352
rect 64980 14288 65044 14352
rect 65060 14288 65124 14352
rect 65140 14288 65204 14352
rect 65220 14288 65284 14352
rect 70740 14288 70804 14352
rect 70820 14288 70884 14352
rect 70900 14288 70964 14352
rect 70980 14288 71044 14352
rect 71060 14288 71124 14352
rect 71140 14288 71204 14352
rect 71220 14288 71284 14352
rect 66852 12684 66916 12748
rect 64092 12548 64156 12612
rect 1740 12176 1804 12240
rect 1820 12176 1884 12240
rect 1900 12176 1964 12240
rect 1980 12176 2044 12240
rect 2060 12176 2124 12240
rect 2140 12176 2204 12240
rect 2220 12176 2284 12240
rect 7740 12176 7804 12240
rect 7820 12176 7884 12240
rect 7900 12176 7964 12240
rect 7980 12176 8044 12240
rect 8060 12176 8124 12240
rect 8140 12176 8204 12240
rect 8220 12176 8284 12240
rect 13740 12176 13804 12240
rect 13820 12176 13884 12240
rect 13900 12176 13964 12240
rect 13980 12176 14044 12240
rect 14060 12176 14124 12240
rect 14140 12176 14204 12240
rect 14220 12176 14284 12240
rect 19740 12176 19804 12240
rect 19820 12176 19884 12240
rect 19900 12176 19964 12240
rect 19980 12176 20044 12240
rect 20060 12176 20124 12240
rect 20140 12176 20204 12240
rect 20220 12176 20284 12240
rect 25740 12176 25804 12240
rect 25820 12176 25884 12240
rect 25900 12176 25964 12240
rect 25980 12176 26044 12240
rect 26060 12176 26124 12240
rect 26140 12176 26204 12240
rect 26220 12176 26284 12240
rect 31740 12176 31804 12240
rect 31820 12176 31884 12240
rect 31900 12176 31964 12240
rect 31980 12176 32044 12240
rect 32060 12176 32124 12240
rect 32140 12176 32204 12240
rect 32220 12176 32284 12240
rect 37740 12176 37804 12240
rect 37820 12176 37884 12240
rect 37900 12176 37964 12240
rect 37980 12176 38044 12240
rect 38060 12176 38124 12240
rect 38140 12176 38204 12240
rect 38220 12176 38284 12240
rect 43740 12176 43804 12240
rect 43820 12176 43884 12240
rect 43900 12176 43964 12240
rect 43980 12176 44044 12240
rect 44060 12176 44124 12240
rect 44140 12176 44204 12240
rect 44220 12176 44284 12240
rect 49740 12176 49804 12240
rect 49820 12176 49884 12240
rect 49900 12176 49964 12240
rect 49980 12176 50044 12240
rect 50060 12176 50124 12240
rect 50140 12176 50204 12240
rect 50220 12176 50284 12240
rect 55740 12176 55804 12240
rect 55820 12176 55884 12240
rect 55900 12176 55964 12240
rect 55980 12176 56044 12240
rect 56060 12176 56124 12240
rect 56140 12176 56204 12240
rect 56220 12176 56284 12240
rect 61740 12176 61804 12240
rect 61820 12176 61884 12240
rect 61900 12176 61964 12240
rect 61980 12176 62044 12240
rect 62060 12176 62124 12240
rect 62140 12176 62204 12240
rect 62220 12176 62284 12240
rect 67740 12176 67804 12240
rect 67820 12176 67884 12240
rect 67900 12176 67964 12240
rect 67980 12176 68044 12240
rect 68060 12176 68124 12240
rect 68140 12176 68204 12240
rect 68220 12176 68284 12240
rect 73740 12176 73804 12240
rect 73820 12176 73884 12240
rect 73900 12176 73964 12240
rect 73980 12176 74044 12240
rect 74060 12176 74124 12240
rect 74140 12176 74204 12240
rect 74220 12176 74284 12240
rect 1740 12096 1804 12160
rect 1820 12096 1884 12160
rect 1900 12096 1964 12160
rect 1980 12096 2044 12160
rect 2060 12096 2124 12160
rect 2140 12096 2204 12160
rect 2220 12096 2284 12160
rect 7740 12096 7804 12160
rect 7820 12096 7884 12160
rect 7900 12096 7964 12160
rect 7980 12096 8044 12160
rect 8060 12096 8124 12160
rect 8140 12096 8204 12160
rect 8220 12096 8284 12160
rect 13740 12096 13804 12160
rect 13820 12096 13884 12160
rect 13900 12096 13964 12160
rect 13980 12096 14044 12160
rect 14060 12096 14124 12160
rect 14140 12096 14204 12160
rect 14220 12096 14284 12160
rect 19740 12096 19804 12160
rect 19820 12096 19884 12160
rect 19900 12096 19964 12160
rect 19980 12096 20044 12160
rect 20060 12096 20124 12160
rect 20140 12096 20204 12160
rect 20220 12096 20284 12160
rect 25740 12096 25804 12160
rect 25820 12096 25884 12160
rect 25900 12096 25964 12160
rect 25980 12096 26044 12160
rect 26060 12096 26124 12160
rect 26140 12096 26204 12160
rect 26220 12096 26284 12160
rect 31740 12096 31804 12160
rect 31820 12096 31884 12160
rect 31900 12096 31964 12160
rect 31980 12096 32044 12160
rect 32060 12096 32124 12160
rect 32140 12096 32204 12160
rect 32220 12096 32284 12160
rect 37740 12096 37804 12160
rect 37820 12096 37884 12160
rect 37900 12096 37964 12160
rect 37980 12096 38044 12160
rect 38060 12096 38124 12160
rect 38140 12096 38204 12160
rect 38220 12096 38284 12160
rect 43740 12096 43804 12160
rect 43820 12096 43884 12160
rect 43900 12096 43964 12160
rect 43980 12096 44044 12160
rect 44060 12096 44124 12160
rect 44140 12096 44204 12160
rect 44220 12096 44284 12160
rect 49740 12096 49804 12160
rect 49820 12096 49884 12160
rect 49900 12096 49964 12160
rect 49980 12096 50044 12160
rect 50060 12096 50124 12160
rect 50140 12096 50204 12160
rect 50220 12096 50284 12160
rect 55740 12096 55804 12160
rect 55820 12096 55884 12160
rect 55900 12096 55964 12160
rect 55980 12096 56044 12160
rect 56060 12096 56124 12160
rect 56140 12096 56204 12160
rect 56220 12096 56284 12160
rect 61740 12096 61804 12160
rect 61820 12096 61884 12160
rect 61900 12096 61964 12160
rect 61980 12096 62044 12160
rect 62060 12096 62124 12160
rect 62140 12096 62204 12160
rect 62220 12096 62284 12160
rect 67740 12096 67804 12160
rect 67820 12096 67884 12160
rect 67900 12096 67964 12160
rect 67980 12096 68044 12160
rect 68060 12096 68124 12160
rect 68140 12096 68204 12160
rect 68220 12096 68284 12160
rect 73740 12096 73804 12160
rect 73820 12096 73884 12160
rect 73900 12096 73964 12160
rect 73980 12096 74044 12160
rect 74060 12096 74124 12160
rect 74140 12096 74204 12160
rect 74220 12096 74284 12160
rect 1740 12016 1804 12080
rect 1820 12016 1884 12080
rect 1900 12016 1964 12080
rect 1980 12016 2044 12080
rect 2060 12016 2124 12080
rect 2140 12016 2204 12080
rect 2220 12016 2284 12080
rect 7740 12016 7804 12080
rect 7820 12016 7884 12080
rect 7900 12016 7964 12080
rect 7980 12016 8044 12080
rect 8060 12016 8124 12080
rect 8140 12016 8204 12080
rect 8220 12016 8284 12080
rect 13740 12016 13804 12080
rect 13820 12016 13884 12080
rect 13900 12016 13964 12080
rect 13980 12016 14044 12080
rect 14060 12016 14124 12080
rect 14140 12016 14204 12080
rect 14220 12016 14284 12080
rect 19740 12016 19804 12080
rect 19820 12016 19884 12080
rect 19900 12016 19964 12080
rect 19980 12016 20044 12080
rect 20060 12016 20124 12080
rect 20140 12016 20204 12080
rect 20220 12016 20284 12080
rect 25740 12016 25804 12080
rect 25820 12016 25884 12080
rect 25900 12016 25964 12080
rect 25980 12016 26044 12080
rect 26060 12016 26124 12080
rect 26140 12016 26204 12080
rect 26220 12016 26284 12080
rect 31740 12016 31804 12080
rect 31820 12016 31884 12080
rect 31900 12016 31964 12080
rect 31980 12016 32044 12080
rect 32060 12016 32124 12080
rect 32140 12016 32204 12080
rect 32220 12016 32284 12080
rect 37740 12016 37804 12080
rect 37820 12016 37884 12080
rect 37900 12016 37964 12080
rect 37980 12016 38044 12080
rect 38060 12016 38124 12080
rect 38140 12016 38204 12080
rect 38220 12016 38284 12080
rect 43740 12016 43804 12080
rect 43820 12016 43884 12080
rect 43900 12016 43964 12080
rect 43980 12016 44044 12080
rect 44060 12016 44124 12080
rect 44140 12016 44204 12080
rect 44220 12016 44284 12080
rect 49740 12016 49804 12080
rect 49820 12016 49884 12080
rect 49900 12016 49964 12080
rect 49980 12016 50044 12080
rect 50060 12016 50124 12080
rect 50140 12016 50204 12080
rect 50220 12016 50284 12080
rect 55740 12016 55804 12080
rect 55820 12016 55884 12080
rect 55900 12016 55964 12080
rect 55980 12016 56044 12080
rect 56060 12016 56124 12080
rect 56140 12016 56204 12080
rect 56220 12016 56284 12080
rect 61740 12016 61804 12080
rect 61820 12016 61884 12080
rect 61900 12016 61964 12080
rect 61980 12016 62044 12080
rect 62060 12016 62124 12080
rect 62140 12016 62204 12080
rect 62220 12016 62284 12080
rect 67740 12016 67804 12080
rect 67820 12016 67884 12080
rect 67900 12016 67964 12080
rect 67980 12016 68044 12080
rect 68060 12016 68124 12080
rect 68140 12016 68204 12080
rect 68220 12016 68284 12080
rect 73740 12016 73804 12080
rect 73820 12016 73884 12080
rect 73900 12016 73964 12080
rect 73980 12016 74044 12080
rect 74060 12016 74124 12080
rect 74140 12016 74204 12080
rect 74220 12016 74284 12080
rect 1740 11936 1804 12000
rect 1820 11936 1884 12000
rect 1900 11936 1964 12000
rect 1980 11936 2044 12000
rect 2060 11936 2124 12000
rect 2140 11936 2204 12000
rect 2220 11936 2284 12000
rect 7740 11936 7804 12000
rect 7820 11936 7884 12000
rect 7900 11936 7964 12000
rect 7980 11936 8044 12000
rect 8060 11936 8124 12000
rect 8140 11936 8204 12000
rect 8220 11936 8284 12000
rect 13740 11936 13804 12000
rect 13820 11936 13884 12000
rect 13900 11936 13964 12000
rect 13980 11936 14044 12000
rect 14060 11936 14124 12000
rect 14140 11936 14204 12000
rect 14220 11936 14284 12000
rect 19740 11936 19804 12000
rect 19820 11936 19884 12000
rect 19900 11936 19964 12000
rect 19980 11936 20044 12000
rect 20060 11936 20124 12000
rect 20140 11936 20204 12000
rect 20220 11936 20284 12000
rect 25740 11936 25804 12000
rect 25820 11936 25884 12000
rect 25900 11936 25964 12000
rect 25980 11936 26044 12000
rect 26060 11936 26124 12000
rect 26140 11936 26204 12000
rect 26220 11936 26284 12000
rect 31740 11936 31804 12000
rect 31820 11936 31884 12000
rect 31900 11936 31964 12000
rect 31980 11936 32044 12000
rect 32060 11936 32124 12000
rect 32140 11936 32204 12000
rect 32220 11936 32284 12000
rect 37740 11936 37804 12000
rect 37820 11936 37884 12000
rect 37900 11936 37964 12000
rect 37980 11936 38044 12000
rect 38060 11936 38124 12000
rect 38140 11936 38204 12000
rect 38220 11936 38284 12000
rect 43740 11936 43804 12000
rect 43820 11936 43884 12000
rect 43900 11936 43964 12000
rect 43980 11936 44044 12000
rect 44060 11936 44124 12000
rect 44140 11936 44204 12000
rect 44220 11936 44284 12000
rect 49740 11936 49804 12000
rect 49820 11936 49884 12000
rect 49900 11936 49964 12000
rect 49980 11936 50044 12000
rect 50060 11936 50124 12000
rect 50140 11936 50204 12000
rect 50220 11936 50284 12000
rect 55740 11936 55804 12000
rect 55820 11936 55884 12000
rect 55900 11936 55964 12000
rect 55980 11936 56044 12000
rect 56060 11936 56124 12000
rect 56140 11936 56204 12000
rect 56220 11936 56284 12000
rect 61740 11936 61804 12000
rect 61820 11936 61884 12000
rect 61900 11936 61964 12000
rect 61980 11936 62044 12000
rect 62060 11936 62124 12000
rect 62140 11936 62204 12000
rect 62220 11936 62284 12000
rect 67740 11936 67804 12000
rect 67820 11936 67884 12000
rect 67900 11936 67964 12000
rect 67980 11936 68044 12000
rect 68060 11936 68124 12000
rect 68140 11936 68204 12000
rect 68220 11936 68284 12000
rect 73740 11936 73804 12000
rect 73820 11936 73884 12000
rect 73900 11936 73964 12000
rect 73980 11936 74044 12000
rect 74060 11936 74124 12000
rect 74140 11936 74204 12000
rect 74220 11936 74284 12000
rect 63540 11792 63604 11796
rect 63540 11736 63554 11792
rect 63554 11736 63604 11792
rect 63540 11732 63604 11736
rect 64276 11732 64340 11796
rect 63356 11596 63420 11660
rect 63908 11596 63972 11660
rect 64092 11052 64156 11116
rect 63356 10704 63420 10708
rect 63356 10648 63406 10704
rect 63406 10648 63420 10704
rect 63356 10644 63420 10648
rect 63908 7652 63972 7716
rect 62988 7516 63052 7580
rect 63356 7244 63420 7308
rect 64092 6972 64156 7036
rect 65564 6700 65628 6764
rect 65748 6564 65812 6628
rect 66484 6292 66548 6356
rect 66852 6156 66916 6220
rect 65932 6020 65996 6084
rect 39988 5748 40052 5812
rect 63172 5748 63236 5812
rect 68508 5612 68572 5676
rect 64276 5068 64340 5132
rect 64460 4932 64524 4996
rect 66668 4796 66732 4860
rect 4740 4528 4804 4592
rect 4820 4528 4884 4592
rect 4900 4528 4964 4592
rect 4980 4528 5044 4592
rect 5060 4528 5124 4592
rect 5140 4528 5204 4592
rect 5220 4528 5284 4592
rect 10740 4528 10804 4592
rect 10820 4528 10884 4592
rect 10900 4528 10964 4592
rect 10980 4528 11044 4592
rect 11060 4528 11124 4592
rect 11140 4528 11204 4592
rect 11220 4528 11284 4592
rect 16740 4528 16804 4592
rect 16820 4528 16884 4592
rect 16900 4528 16964 4592
rect 16980 4528 17044 4592
rect 17060 4528 17124 4592
rect 17140 4528 17204 4592
rect 17220 4528 17284 4592
rect 22740 4528 22804 4592
rect 22820 4528 22884 4592
rect 22900 4528 22964 4592
rect 22980 4528 23044 4592
rect 23060 4528 23124 4592
rect 23140 4528 23204 4592
rect 23220 4528 23284 4592
rect 28740 4528 28804 4592
rect 28820 4528 28884 4592
rect 28900 4528 28964 4592
rect 28980 4528 29044 4592
rect 29060 4528 29124 4592
rect 29140 4528 29204 4592
rect 29220 4528 29284 4592
rect 34740 4528 34804 4592
rect 34820 4528 34884 4592
rect 34900 4528 34964 4592
rect 34980 4528 35044 4592
rect 35060 4528 35124 4592
rect 35140 4528 35204 4592
rect 35220 4528 35284 4592
rect 40740 4528 40804 4592
rect 40820 4528 40884 4592
rect 40900 4528 40964 4592
rect 40980 4528 41044 4592
rect 41060 4528 41124 4592
rect 41140 4528 41204 4592
rect 41220 4528 41284 4592
rect 46740 4528 46804 4592
rect 46820 4528 46884 4592
rect 46900 4528 46964 4592
rect 46980 4528 47044 4592
rect 47060 4528 47124 4592
rect 47140 4528 47204 4592
rect 47220 4528 47284 4592
rect 52740 4528 52804 4592
rect 52820 4528 52884 4592
rect 52900 4528 52964 4592
rect 52980 4528 53044 4592
rect 53060 4528 53124 4592
rect 53140 4528 53204 4592
rect 53220 4528 53284 4592
rect 58740 4528 58804 4592
rect 58820 4528 58884 4592
rect 58900 4528 58964 4592
rect 58980 4528 59044 4592
rect 59060 4528 59124 4592
rect 59140 4528 59204 4592
rect 59220 4528 59284 4592
rect 64740 4528 64804 4592
rect 64820 4528 64884 4592
rect 64900 4528 64964 4592
rect 64980 4528 65044 4592
rect 65060 4528 65124 4592
rect 65140 4528 65204 4592
rect 65220 4528 65284 4592
rect 70740 4528 70804 4592
rect 70820 4528 70884 4592
rect 70900 4528 70964 4592
rect 70980 4528 71044 4592
rect 71060 4528 71124 4592
rect 71140 4528 71204 4592
rect 71220 4528 71284 4592
rect 4740 4448 4804 4512
rect 4820 4448 4884 4512
rect 4900 4448 4964 4512
rect 4980 4448 5044 4512
rect 5060 4448 5124 4512
rect 5140 4448 5204 4512
rect 5220 4448 5284 4512
rect 10740 4448 10804 4512
rect 10820 4448 10884 4512
rect 10900 4448 10964 4512
rect 10980 4448 11044 4512
rect 11060 4448 11124 4512
rect 11140 4448 11204 4512
rect 11220 4448 11284 4512
rect 16740 4448 16804 4512
rect 16820 4448 16884 4512
rect 16900 4448 16964 4512
rect 16980 4448 17044 4512
rect 17060 4448 17124 4512
rect 17140 4448 17204 4512
rect 17220 4448 17284 4512
rect 22740 4448 22804 4512
rect 22820 4448 22884 4512
rect 22900 4448 22964 4512
rect 22980 4448 23044 4512
rect 23060 4448 23124 4512
rect 23140 4448 23204 4512
rect 23220 4448 23284 4512
rect 28740 4448 28804 4512
rect 28820 4448 28884 4512
rect 28900 4448 28964 4512
rect 28980 4448 29044 4512
rect 29060 4448 29124 4512
rect 29140 4448 29204 4512
rect 29220 4448 29284 4512
rect 34740 4448 34804 4512
rect 34820 4448 34884 4512
rect 34900 4448 34964 4512
rect 34980 4448 35044 4512
rect 35060 4448 35124 4512
rect 35140 4448 35204 4512
rect 35220 4448 35284 4512
rect 40740 4448 40804 4512
rect 40820 4448 40884 4512
rect 40900 4448 40964 4512
rect 40980 4448 41044 4512
rect 41060 4448 41124 4512
rect 41140 4448 41204 4512
rect 41220 4448 41284 4512
rect 46740 4448 46804 4512
rect 46820 4448 46884 4512
rect 46900 4448 46964 4512
rect 46980 4448 47044 4512
rect 47060 4448 47124 4512
rect 47140 4448 47204 4512
rect 47220 4448 47284 4512
rect 52740 4448 52804 4512
rect 52820 4448 52884 4512
rect 52900 4448 52964 4512
rect 52980 4448 53044 4512
rect 53060 4448 53124 4512
rect 53140 4448 53204 4512
rect 53220 4448 53284 4512
rect 58740 4448 58804 4512
rect 58820 4448 58884 4512
rect 58900 4448 58964 4512
rect 58980 4448 59044 4512
rect 59060 4448 59124 4512
rect 59140 4448 59204 4512
rect 59220 4448 59284 4512
rect 64740 4448 64804 4512
rect 64820 4448 64884 4512
rect 64900 4448 64964 4512
rect 64980 4448 65044 4512
rect 65060 4448 65124 4512
rect 65140 4448 65204 4512
rect 65220 4448 65284 4512
rect 70740 4448 70804 4512
rect 70820 4448 70884 4512
rect 70900 4448 70964 4512
rect 70980 4448 71044 4512
rect 71060 4448 71124 4512
rect 71140 4448 71204 4512
rect 71220 4448 71284 4512
rect 4740 4368 4804 4432
rect 4820 4368 4884 4432
rect 4900 4368 4964 4432
rect 4980 4368 5044 4432
rect 5060 4368 5124 4432
rect 5140 4368 5204 4432
rect 5220 4368 5284 4432
rect 10740 4368 10804 4432
rect 10820 4368 10884 4432
rect 10900 4368 10964 4432
rect 10980 4368 11044 4432
rect 11060 4368 11124 4432
rect 11140 4368 11204 4432
rect 11220 4368 11284 4432
rect 16740 4368 16804 4432
rect 16820 4368 16884 4432
rect 16900 4368 16964 4432
rect 16980 4368 17044 4432
rect 17060 4368 17124 4432
rect 17140 4368 17204 4432
rect 17220 4368 17284 4432
rect 22740 4368 22804 4432
rect 22820 4368 22884 4432
rect 22900 4368 22964 4432
rect 22980 4368 23044 4432
rect 23060 4368 23124 4432
rect 23140 4368 23204 4432
rect 23220 4368 23284 4432
rect 28740 4368 28804 4432
rect 28820 4368 28884 4432
rect 28900 4368 28964 4432
rect 28980 4368 29044 4432
rect 29060 4368 29124 4432
rect 29140 4368 29204 4432
rect 29220 4368 29284 4432
rect 34740 4368 34804 4432
rect 34820 4368 34884 4432
rect 34900 4368 34964 4432
rect 34980 4368 35044 4432
rect 35060 4368 35124 4432
rect 35140 4368 35204 4432
rect 35220 4368 35284 4432
rect 40740 4368 40804 4432
rect 40820 4368 40884 4432
rect 40900 4368 40964 4432
rect 40980 4368 41044 4432
rect 41060 4368 41124 4432
rect 41140 4368 41204 4432
rect 41220 4368 41284 4432
rect 46740 4368 46804 4432
rect 46820 4368 46884 4432
rect 46900 4368 46964 4432
rect 46980 4368 47044 4432
rect 47060 4368 47124 4432
rect 47140 4368 47204 4432
rect 47220 4368 47284 4432
rect 52740 4368 52804 4432
rect 52820 4368 52884 4432
rect 52900 4368 52964 4432
rect 52980 4368 53044 4432
rect 53060 4368 53124 4432
rect 53140 4368 53204 4432
rect 53220 4368 53284 4432
rect 58740 4368 58804 4432
rect 58820 4368 58884 4432
rect 58900 4368 58964 4432
rect 58980 4368 59044 4432
rect 59060 4368 59124 4432
rect 59140 4368 59204 4432
rect 59220 4368 59284 4432
rect 64740 4368 64804 4432
rect 64820 4368 64884 4432
rect 64900 4368 64964 4432
rect 64980 4368 65044 4432
rect 65060 4368 65124 4432
rect 65140 4368 65204 4432
rect 65220 4368 65284 4432
rect 70740 4368 70804 4432
rect 70820 4368 70884 4432
rect 70900 4368 70964 4432
rect 70980 4368 71044 4432
rect 71060 4368 71124 4432
rect 71140 4368 71204 4432
rect 71220 4368 71284 4432
rect 4740 4288 4804 4352
rect 4820 4288 4884 4352
rect 4900 4288 4964 4352
rect 4980 4288 5044 4352
rect 5060 4288 5124 4352
rect 5140 4288 5204 4352
rect 5220 4288 5284 4352
rect 10740 4288 10804 4352
rect 10820 4288 10884 4352
rect 10900 4288 10964 4352
rect 10980 4288 11044 4352
rect 11060 4288 11124 4352
rect 11140 4288 11204 4352
rect 11220 4288 11284 4352
rect 16740 4288 16804 4352
rect 16820 4288 16884 4352
rect 16900 4288 16964 4352
rect 16980 4288 17044 4352
rect 17060 4288 17124 4352
rect 17140 4288 17204 4352
rect 17220 4288 17284 4352
rect 22740 4288 22804 4352
rect 22820 4288 22884 4352
rect 22900 4288 22964 4352
rect 22980 4288 23044 4352
rect 23060 4288 23124 4352
rect 23140 4288 23204 4352
rect 23220 4288 23284 4352
rect 28740 4288 28804 4352
rect 28820 4288 28884 4352
rect 28900 4288 28964 4352
rect 28980 4288 29044 4352
rect 29060 4288 29124 4352
rect 29140 4288 29204 4352
rect 29220 4288 29284 4352
rect 34740 4288 34804 4352
rect 34820 4288 34884 4352
rect 34900 4288 34964 4352
rect 34980 4288 35044 4352
rect 35060 4288 35124 4352
rect 35140 4288 35204 4352
rect 35220 4288 35284 4352
rect 40740 4288 40804 4352
rect 40820 4288 40884 4352
rect 40900 4288 40964 4352
rect 40980 4288 41044 4352
rect 41060 4288 41124 4352
rect 41140 4288 41204 4352
rect 41220 4288 41284 4352
rect 46740 4288 46804 4352
rect 46820 4288 46884 4352
rect 46900 4288 46964 4352
rect 46980 4288 47044 4352
rect 47060 4288 47124 4352
rect 47140 4288 47204 4352
rect 47220 4288 47284 4352
rect 52740 4288 52804 4352
rect 52820 4288 52884 4352
rect 52900 4288 52964 4352
rect 52980 4288 53044 4352
rect 53060 4288 53124 4352
rect 53140 4288 53204 4352
rect 53220 4288 53284 4352
rect 58740 4288 58804 4352
rect 58820 4288 58884 4352
rect 58900 4288 58964 4352
rect 58980 4288 59044 4352
rect 59060 4288 59124 4352
rect 59140 4288 59204 4352
rect 59220 4288 59284 4352
rect 64740 4288 64804 4352
rect 64820 4288 64884 4352
rect 64900 4288 64964 4352
rect 64980 4288 65044 4352
rect 65060 4288 65124 4352
rect 65140 4288 65204 4352
rect 65220 4288 65284 4352
rect 70740 4288 70804 4352
rect 70820 4288 70884 4352
rect 70900 4288 70964 4352
rect 70980 4288 71044 4352
rect 71060 4288 71124 4352
rect 71140 4288 71204 4352
rect 71220 4288 71284 4352
rect 63724 3980 63788 4044
rect 39988 3300 40052 3364
rect 66300 3300 66364 3364
rect 1740 2176 1804 2240
rect 1820 2236 1884 2240
rect 1900 2236 1964 2240
rect 1980 2236 2044 2240
rect 2060 2236 2124 2240
rect 2140 2236 2204 2240
rect 1820 2180 1864 2236
rect 1864 2180 1884 2236
rect 1900 2180 1920 2236
rect 1920 2180 1944 2236
rect 1944 2180 1964 2236
rect 1980 2180 2000 2236
rect 2000 2180 2024 2236
rect 2024 2180 2044 2236
rect 2060 2180 2080 2236
rect 2080 2180 2104 2236
rect 2104 2180 2124 2236
rect 2140 2180 2160 2236
rect 2160 2180 2204 2236
rect 1820 2176 1884 2180
rect 1900 2176 1964 2180
rect 1980 2176 2044 2180
rect 2060 2176 2124 2180
rect 2140 2176 2204 2180
rect 2220 2176 2284 2240
rect 7740 2176 7804 2240
rect 7820 2176 7884 2240
rect 7900 2176 7964 2240
rect 7980 2176 8044 2240
rect 8060 2176 8124 2240
rect 8140 2176 8204 2240
rect 8220 2176 8284 2240
rect 13740 2176 13804 2240
rect 13820 2176 13884 2240
rect 13900 2176 13964 2240
rect 13980 2176 14044 2240
rect 14060 2176 14124 2240
rect 14140 2176 14204 2240
rect 14220 2176 14284 2240
rect 19740 2176 19804 2240
rect 19820 2176 19884 2240
rect 19900 2176 19964 2240
rect 19980 2176 20044 2240
rect 20060 2176 20124 2240
rect 20140 2176 20204 2240
rect 20220 2176 20284 2240
rect 25740 2176 25804 2240
rect 25820 2176 25884 2240
rect 25900 2176 25964 2240
rect 25980 2176 26044 2240
rect 26060 2176 26124 2240
rect 26140 2176 26204 2240
rect 26220 2176 26284 2240
rect 31740 2176 31804 2240
rect 31820 2236 31884 2240
rect 31900 2236 31964 2240
rect 31980 2236 32044 2240
rect 32060 2236 32124 2240
rect 32140 2236 32204 2240
rect 31820 2180 31864 2236
rect 31864 2180 31884 2236
rect 31900 2180 31920 2236
rect 31920 2180 31944 2236
rect 31944 2180 31964 2236
rect 31980 2180 32000 2236
rect 32000 2180 32024 2236
rect 32024 2180 32044 2236
rect 32060 2180 32080 2236
rect 32080 2180 32104 2236
rect 32104 2180 32124 2236
rect 32140 2180 32160 2236
rect 32160 2180 32204 2236
rect 31820 2176 31884 2180
rect 31900 2176 31964 2180
rect 31980 2176 32044 2180
rect 32060 2176 32124 2180
rect 32140 2176 32204 2180
rect 32220 2176 32284 2240
rect 37740 2176 37804 2240
rect 37820 2176 37884 2240
rect 37900 2176 37964 2240
rect 37980 2176 38044 2240
rect 38060 2176 38124 2240
rect 38140 2176 38204 2240
rect 38220 2176 38284 2240
rect 43740 2176 43804 2240
rect 43820 2176 43884 2240
rect 43900 2176 43964 2240
rect 43980 2176 44044 2240
rect 44060 2176 44124 2240
rect 44140 2176 44204 2240
rect 44220 2176 44284 2240
rect 49740 2176 49804 2240
rect 49820 2176 49884 2240
rect 49900 2176 49964 2240
rect 49980 2176 50044 2240
rect 50060 2176 50124 2240
rect 50140 2176 50204 2240
rect 50220 2176 50284 2240
rect 55740 2176 55804 2240
rect 55820 2176 55884 2240
rect 55900 2176 55964 2240
rect 55980 2176 56044 2240
rect 56060 2176 56124 2240
rect 56140 2176 56204 2240
rect 56220 2176 56284 2240
rect 61740 2176 61804 2240
rect 61820 2236 61884 2240
rect 61900 2236 61964 2240
rect 61980 2236 62044 2240
rect 62060 2236 62124 2240
rect 62140 2236 62204 2240
rect 61820 2180 61864 2236
rect 61864 2180 61884 2236
rect 61900 2180 61920 2236
rect 61920 2180 61944 2236
rect 61944 2180 61964 2236
rect 61980 2180 62000 2236
rect 62000 2180 62024 2236
rect 62024 2180 62044 2236
rect 62060 2180 62080 2236
rect 62080 2180 62104 2236
rect 62104 2180 62124 2236
rect 62140 2180 62160 2236
rect 62160 2180 62204 2236
rect 61820 2176 61884 2180
rect 61900 2176 61964 2180
rect 61980 2176 62044 2180
rect 62060 2176 62124 2180
rect 62140 2176 62204 2180
rect 62220 2176 62284 2240
rect 67740 2176 67804 2240
rect 67820 2176 67884 2240
rect 67900 2176 67964 2240
rect 67980 2176 68044 2240
rect 68060 2176 68124 2240
rect 68140 2176 68204 2240
rect 68220 2176 68284 2240
rect 73740 2176 73804 2240
rect 73820 2176 73884 2240
rect 73900 2176 73964 2240
rect 73980 2176 74044 2240
rect 74060 2176 74124 2240
rect 74140 2176 74204 2240
rect 74220 2176 74284 2240
rect 1740 2096 1804 2160
rect 1820 2156 1884 2160
rect 1900 2156 1964 2160
rect 1980 2156 2044 2160
rect 2060 2156 2124 2160
rect 2140 2156 2204 2160
rect 1820 2100 1864 2156
rect 1864 2100 1884 2156
rect 1900 2100 1920 2156
rect 1920 2100 1944 2156
rect 1944 2100 1964 2156
rect 1980 2100 2000 2156
rect 2000 2100 2024 2156
rect 2024 2100 2044 2156
rect 2060 2100 2080 2156
rect 2080 2100 2104 2156
rect 2104 2100 2124 2156
rect 2140 2100 2160 2156
rect 2160 2100 2204 2156
rect 1820 2096 1884 2100
rect 1900 2096 1964 2100
rect 1980 2096 2044 2100
rect 2060 2096 2124 2100
rect 2140 2096 2204 2100
rect 2220 2096 2284 2160
rect 7740 2096 7804 2160
rect 7820 2096 7884 2160
rect 7900 2096 7964 2160
rect 7980 2096 8044 2160
rect 8060 2096 8124 2160
rect 8140 2096 8204 2160
rect 8220 2096 8284 2160
rect 13740 2096 13804 2160
rect 13820 2096 13884 2160
rect 13900 2096 13964 2160
rect 13980 2096 14044 2160
rect 14060 2096 14124 2160
rect 14140 2096 14204 2160
rect 14220 2096 14284 2160
rect 19740 2096 19804 2160
rect 19820 2096 19884 2160
rect 19900 2096 19964 2160
rect 19980 2096 20044 2160
rect 20060 2096 20124 2160
rect 20140 2096 20204 2160
rect 20220 2096 20284 2160
rect 25740 2096 25804 2160
rect 25820 2096 25884 2160
rect 25900 2096 25964 2160
rect 25980 2096 26044 2160
rect 26060 2096 26124 2160
rect 26140 2096 26204 2160
rect 26220 2096 26284 2160
rect 31740 2096 31804 2160
rect 31820 2156 31884 2160
rect 31900 2156 31964 2160
rect 31980 2156 32044 2160
rect 32060 2156 32124 2160
rect 32140 2156 32204 2160
rect 31820 2100 31864 2156
rect 31864 2100 31884 2156
rect 31900 2100 31920 2156
rect 31920 2100 31944 2156
rect 31944 2100 31964 2156
rect 31980 2100 32000 2156
rect 32000 2100 32024 2156
rect 32024 2100 32044 2156
rect 32060 2100 32080 2156
rect 32080 2100 32104 2156
rect 32104 2100 32124 2156
rect 32140 2100 32160 2156
rect 32160 2100 32204 2156
rect 31820 2096 31884 2100
rect 31900 2096 31964 2100
rect 31980 2096 32044 2100
rect 32060 2096 32124 2100
rect 32140 2096 32204 2100
rect 32220 2096 32284 2160
rect 37740 2096 37804 2160
rect 37820 2096 37884 2160
rect 37900 2096 37964 2160
rect 37980 2096 38044 2160
rect 38060 2096 38124 2160
rect 38140 2096 38204 2160
rect 38220 2096 38284 2160
rect 43740 2096 43804 2160
rect 43820 2096 43884 2160
rect 43900 2096 43964 2160
rect 43980 2096 44044 2160
rect 44060 2096 44124 2160
rect 44140 2096 44204 2160
rect 44220 2096 44284 2160
rect 49740 2096 49804 2160
rect 49820 2096 49884 2160
rect 49900 2096 49964 2160
rect 49980 2096 50044 2160
rect 50060 2096 50124 2160
rect 50140 2096 50204 2160
rect 50220 2096 50284 2160
rect 55740 2096 55804 2160
rect 55820 2096 55884 2160
rect 55900 2096 55964 2160
rect 55980 2096 56044 2160
rect 56060 2096 56124 2160
rect 56140 2096 56204 2160
rect 56220 2096 56284 2160
rect 61740 2096 61804 2160
rect 61820 2156 61884 2160
rect 61900 2156 61964 2160
rect 61980 2156 62044 2160
rect 62060 2156 62124 2160
rect 62140 2156 62204 2160
rect 61820 2100 61864 2156
rect 61864 2100 61884 2156
rect 61900 2100 61920 2156
rect 61920 2100 61944 2156
rect 61944 2100 61964 2156
rect 61980 2100 62000 2156
rect 62000 2100 62024 2156
rect 62024 2100 62044 2156
rect 62060 2100 62080 2156
rect 62080 2100 62104 2156
rect 62104 2100 62124 2156
rect 62140 2100 62160 2156
rect 62160 2100 62204 2156
rect 61820 2096 61884 2100
rect 61900 2096 61964 2100
rect 61980 2096 62044 2100
rect 62060 2096 62124 2100
rect 62140 2096 62204 2100
rect 62220 2096 62284 2160
rect 67740 2096 67804 2160
rect 67820 2096 67884 2160
rect 67900 2096 67964 2160
rect 67980 2096 68044 2160
rect 68060 2096 68124 2160
rect 68140 2096 68204 2160
rect 68220 2096 68284 2160
rect 73740 2096 73804 2160
rect 73820 2096 73884 2160
rect 73900 2096 73964 2160
rect 73980 2096 74044 2160
rect 74060 2096 74124 2160
rect 74140 2096 74204 2160
rect 74220 2096 74284 2160
rect 1740 2016 1804 2080
rect 1820 2076 1884 2080
rect 1900 2076 1964 2080
rect 1980 2076 2044 2080
rect 2060 2076 2124 2080
rect 2140 2076 2204 2080
rect 1820 2020 1864 2076
rect 1864 2020 1884 2076
rect 1900 2020 1920 2076
rect 1920 2020 1944 2076
rect 1944 2020 1964 2076
rect 1980 2020 2000 2076
rect 2000 2020 2024 2076
rect 2024 2020 2044 2076
rect 2060 2020 2080 2076
rect 2080 2020 2104 2076
rect 2104 2020 2124 2076
rect 2140 2020 2160 2076
rect 2160 2020 2204 2076
rect 1820 2016 1884 2020
rect 1900 2016 1964 2020
rect 1980 2016 2044 2020
rect 2060 2016 2124 2020
rect 2140 2016 2204 2020
rect 2220 2016 2284 2080
rect 7740 2016 7804 2080
rect 7820 2016 7884 2080
rect 7900 2016 7964 2080
rect 7980 2016 8044 2080
rect 8060 2016 8124 2080
rect 8140 2016 8204 2080
rect 8220 2016 8284 2080
rect 13740 2016 13804 2080
rect 13820 2016 13884 2080
rect 13900 2016 13964 2080
rect 13980 2016 14044 2080
rect 14060 2016 14124 2080
rect 14140 2016 14204 2080
rect 14220 2016 14284 2080
rect 19740 2016 19804 2080
rect 19820 2016 19884 2080
rect 19900 2016 19964 2080
rect 19980 2016 20044 2080
rect 20060 2016 20124 2080
rect 20140 2016 20204 2080
rect 20220 2016 20284 2080
rect 25740 2016 25804 2080
rect 25820 2016 25884 2080
rect 25900 2016 25964 2080
rect 25980 2016 26044 2080
rect 26060 2016 26124 2080
rect 26140 2016 26204 2080
rect 26220 2016 26284 2080
rect 31740 2016 31804 2080
rect 31820 2076 31884 2080
rect 31900 2076 31964 2080
rect 31980 2076 32044 2080
rect 32060 2076 32124 2080
rect 32140 2076 32204 2080
rect 31820 2020 31864 2076
rect 31864 2020 31884 2076
rect 31900 2020 31920 2076
rect 31920 2020 31944 2076
rect 31944 2020 31964 2076
rect 31980 2020 32000 2076
rect 32000 2020 32024 2076
rect 32024 2020 32044 2076
rect 32060 2020 32080 2076
rect 32080 2020 32104 2076
rect 32104 2020 32124 2076
rect 32140 2020 32160 2076
rect 32160 2020 32204 2076
rect 31820 2016 31884 2020
rect 31900 2016 31964 2020
rect 31980 2016 32044 2020
rect 32060 2016 32124 2020
rect 32140 2016 32204 2020
rect 32220 2016 32284 2080
rect 37740 2016 37804 2080
rect 37820 2016 37884 2080
rect 37900 2016 37964 2080
rect 37980 2016 38044 2080
rect 38060 2016 38124 2080
rect 38140 2016 38204 2080
rect 38220 2016 38284 2080
rect 43740 2016 43804 2080
rect 43820 2016 43884 2080
rect 43900 2016 43964 2080
rect 43980 2016 44044 2080
rect 44060 2016 44124 2080
rect 44140 2016 44204 2080
rect 44220 2016 44284 2080
rect 49740 2016 49804 2080
rect 49820 2016 49884 2080
rect 49900 2016 49964 2080
rect 49980 2016 50044 2080
rect 50060 2016 50124 2080
rect 50140 2016 50204 2080
rect 50220 2016 50284 2080
rect 55740 2016 55804 2080
rect 55820 2016 55884 2080
rect 55900 2016 55964 2080
rect 55980 2016 56044 2080
rect 56060 2016 56124 2080
rect 56140 2016 56204 2080
rect 56220 2016 56284 2080
rect 61740 2016 61804 2080
rect 61820 2076 61884 2080
rect 61900 2076 61964 2080
rect 61980 2076 62044 2080
rect 62060 2076 62124 2080
rect 62140 2076 62204 2080
rect 61820 2020 61864 2076
rect 61864 2020 61884 2076
rect 61900 2020 61920 2076
rect 61920 2020 61944 2076
rect 61944 2020 61964 2076
rect 61980 2020 62000 2076
rect 62000 2020 62024 2076
rect 62024 2020 62044 2076
rect 62060 2020 62080 2076
rect 62080 2020 62104 2076
rect 62104 2020 62124 2076
rect 62140 2020 62160 2076
rect 62160 2020 62204 2076
rect 61820 2016 61884 2020
rect 61900 2016 61964 2020
rect 61980 2016 62044 2020
rect 62060 2016 62124 2020
rect 62140 2016 62204 2020
rect 62220 2016 62284 2080
rect 67740 2016 67804 2080
rect 67820 2016 67884 2080
rect 67900 2016 67964 2080
rect 67980 2016 68044 2080
rect 68060 2016 68124 2080
rect 68140 2016 68204 2080
rect 68220 2016 68284 2080
rect 73740 2016 73804 2080
rect 73820 2016 73884 2080
rect 73900 2016 73964 2080
rect 73980 2016 74044 2080
rect 74060 2016 74124 2080
rect 74140 2016 74204 2080
rect 74220 2016 74284 2080
rect 1740 1936 1804 2000
rect 1820 1996 1884 2000
rect 1900 1996 1964 2000
rect 1980 1996 2044 2000
rect 2060 1996 2124 2000
rect 2140 1996 2204 2000
rect 1820 1940 1864 1996
rect 1864 1940 1884 1996
rect 1900 1940 1920 1996
rect 1920 1940 1944 1996
rect 1944 1940 1964 1996
rect 1980 1940 2000 1996
rect 2000 1940 2024 1996
rect 2024 1940 2044 1996
rect 2060 1940 2080 1996
rect 2080 1940 2104 1996
rect 2104 1940 2124 1996
rect 2140 1940 2160 1996
rect 2160 1940 2204 1996
rect 1820 1936 1884 1940
rect 1900 1936 1964 1940
rect 1980 1936 2044 1940
rect 2060 1936 2124 1940
rect 2140 1936 2204 1940
rect 2220 1936 2284 2000
rect 7740 1936 7804 2000
rect 7820 1936 7884 2000
rect 7900 1936 7964 2000
rect 7980 1936 8044 2000
rect 8060 1936 8124 2000
rect 8140 1936 8204 2000
rect 8220 1936 8284 2000
rect 13740 1936 13804 2000
rect 13820 1936 13884 2000
rect 13900 1936 13964 2000
rect 13980 1936 14044 2000
rect 14060 1936 14124 2000
rect 14140 1936 14204 2000
rect 14220 1936 14284 2000
rect 19740 1936 19804 2000
rect 19820 1936 19884 2000
rect 19900 1936 19964 2000
rect 19980 1936 20044 2000
rect 20060 1936 20124 2000
rect 20140 1936 20204 2000
rect 20220 1936 20284 2000
rect 25740 1936 25804 2000
rect 25820 1936 25884 2000
rect 25900 1936 25964 2000
rect 25980 1936 26044 2000
rect 26060 1936 26124 2000
rect 26140 1936 26204 2000
rect 26220 1936 26284 2000
rect 31740 1936 31804 2000
rect 31820 1996 31884 2000
rect 31900 1996 31964 2000
rect 31980 1996 32044 2000
rect 32060 1996 32124 2000
rect 32140 1996 32204 2000
rect 31820 1940 31864 1996
rect 31864 1940 31884 1996
rect 31900 1940 31920 1996
rect 31920 1940 31944 1996
rect 31944 1940 31964 1996
rect 31980 1940 32000 1996
rect 32000 1940 32024 1996
rect 32024 1940 32044 1996
rect 32060 1940 32080 1996
rect 32080 1940 32104 1996
rect 32104 1940 32124 1996
rect 32140 1940 32160 1996
rect 32160 1940 32204 1996
rect 31820 1936 31884 1940
rect 31900 1936 31964 1940
rect 31980 1936 32044 1940
rect 32060 1936 32124 1940
rect 32140 1936 32204 1940
rect 32220 1936 32284 2000
rect 37740 1936 37804 2000
rect 37820 1936 37884 2000
rect 37900 1936 37964 2000
rect 37980 1936 38044 2000
rect 38060 1936 38124 2000
rect 38140 1936 38204 2000
rect 38220 1936 38284 2000
rect 43740 1936 43804 2000
rect 43820 1936 43884 2000
rect 43900 1936 43964 2000
rect 43980 1936 44044 2000
rect 44060 1936 44124 2000
rect 44140 1936 44204 2000
rect 44220 1936 44284 2000
rect 49740 1936 49804 2000
rect 49820 1936 49884 2000
rect 49900 1936 49964 2000
rect 49980 1936 50044 2000
rect 50060 1936 50124 2000
rect 50140 1936 50204 2000
rect 50220 1936 50284 2000
rect 55740 1936 55804 2000
rect 55820 1936 55884 2000
rect 55900 1936 55964 2000
rect 55980 1936 56044 2000
rect 56060 1936 56124 2000
rect 56140 1936 56204 2000
rect 56220 1936 56284 2000
rect 61740 1936 61804 2000
rect 61820 1996 61884 2000
rect 61900 1996 61964 2000
rect 61980 1996 62044 2000
rect 62060 1996 62124 2000
rect 62140 1996 62204 2000
rect 61820 1940 61864 1996
rect 61864 1940 61884 1996
rect 61900 1940 61920 1996
rect 61920 1940 61944 1996
rect 61944 1940 61964 1996
rect 61980 1940 62000 1996
rect 62000 1940 62024 1996
rect 62024 1940 62044 1996
rect 62060 1940 62080 1996
rect 62080 1940 62104 1996
rect 62104 1940 62124 1996
rect 62140 1940 62160 1996
rect 62160 1940 62204 1996
rect 61820 1936 61884 1940
rect 61900 1936 61964 1940
rect 61980 1936 62044 1940
rect 62060 1936 62124 1940
rect 62140 1936 62204 1940
rect 62220 1936 62284 2000
rect 67740 1936 67804 2000
rect 67820 1936 67884 2000
rect 67900 1936 67964 2000
rect 67980 1936 68044 2000
rect 68060 1936 68124 2000
rect 68140 1936 68204 2000
rect 68220 1936 68284 2000
rect 73740 1936 73804 2000
rect 73820 1936 73884 2000
rect 73900 1936 73964 2000
rect 73980 1936 74044 2000
rect 74060 1936 74124 2000
rect 74140 1936 74204 2000
rect 74220 1936 74284 2000
<< metal4 >>
rect 1702 82240 2322 87000
rect 1702 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82176 2220 82240
rect 2284 82176 2322 82240
rect 1702 82160 2322 82176
rect 1702 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82096 2220 82160
rect 2284 82096 2322 82160
rect 1702 82080 2322 82096
rect 1702 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82016 2220 82080
rect 2284 82016 2322 82080
rect 1702 82000 2322 82016
rect 1702 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81936 2220 82000
rect 2284 81936 2322 82000
rect 1702 72240 2322 81936
rect 1702 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72176 2220 72240
rect 2284 72176 2322 72240
rect 1702 72160 2322 72176
rect 1702 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72096 2220 72160
rect 2284 72096 2322 72160
rect 1702 72080 2322 72096
rect 1702 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72016 2220 72080
rect 2284 72016 2322 72080
rect 1702 72000 2322 72016
rect 1702 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71936 2220 72000
rect 2284 71936 2322 72000
rect 1702 62240 2322 71936
rect 1702 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62176 2220 62240
rect 2284 62176 2322 62240
rect 1702 62160 2322 62176
rect 1702 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62096 2220 62160
rect 2284 62096 2322 62160
rect 1702 62080 2322 62096
rect 1702 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62016 2220 62080
rect 2284 62016 2322 62080
rect 1702 62000 2322 62016
rect 1702 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61936 2220 62000
rect 2284 61936 2322 62000
rect 1702 52240 2322 61936
rect 1702 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52176 2220 52240
rect 2284 52176 2322 52240
rect 1702 52160 2322 52176
rect 1702 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52096 2220 52160
rect 2284 52096 2322 52160
rect 1702 52080 2322 52096
rect 1702 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52016 2220 52080
rect 2284 52016 2322 52080
rect 1702 52000 2322 52016
rect 1702 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51936 2220 52000
rect 2284 51936 2322 52000
rect 1702 42240 2322 51936
rect 1702 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42176 2220 42240
rect 2284 42176 2322 42240
rect 1702 42160 2322 42176
rect 1702 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42096 2220 42160
rect 2284 42096 2322 42160
rect 1702 42080 2322 42096
rect 1702 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42016 2220 42080
rect 2284 42016 2322 42080
rect 1702 42000 2322 42016
rect 1702 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41936 2220 42000
rect 2284 41936 2322 42000
rect 1702 32240 2322 41936
rect 1702 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32176 2220 32240
rect 2284 32176 2322 32240
rect 1702 32160 2322 32176
rect 1702 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32096 2220 32160
rect 2284 32096 2322 32160
rect 1702 32080 2322 32096
rect 1702 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32016 2220 32080
rect 2284 32016 2322 32080
rect 1702 32000 2322 32016
rect 1702 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31936 2220 32000
rect 2284 31936 2322 32000
rect 1702 22240 2322 31936
rect 1702 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22176 2220 22240
rect 2284 22176 2322 22240
rect 1702 22160 2322 22176
rect 1702 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22096 2220 22160
rect 2284 22096 2322 22160
rect 1702 22080 2322 22096
rect 1702 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22016 2220 22080
rect 2284 22016 2322 22080
rect 1702 22000 2322 22016
rect 1702 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21936 2220 22000
rect 2284 21936 2322 22000
rect 1702 12240 2322 21936
rect 1702 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12176 2220 12240
rect 2284 12176 2322 12240
rect 1702 12160 2322 12176
rect 1702 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12096 2220 12160
rect 2284 12096 2322 12160
rect 1702 12080 2322 12096
rect 1702 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12016 2220 12080
rect 2284 12016 2322 12080
rect 1702 12000 2322 12016
rect 1702 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2220 12000
rect 2284 11936 2322 12000
rect 1702 2240 2322 11936
rect 1702 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2176 1900 2240
rect 1964 2176 1980 2240
rect 2044 2176 2060 2240
rect 2124 2176 2140 2240
rect 2204 2176 2220 2240
rect 2284 2176 2322 2240
rect 1702 2160 2322 2176
rect 1702 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2096 1900 2160
rect 1964 2096 1980 2160
rect 2044 2096 2060 2160
rect 2124 2096 2140 2160
rect 2204 2096 2220 2160
rect 2284 2096 2322 2160
rect 1702 2080 2322 2096
rect 1702 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2016 1900 2080
rect 1964 2016 1980 2080
rect 2044 2016 2060 2080
rect 2124 2016 2140 2080
rect 2204 2016 2220 2080
rect 2284 2016 2322 2080
rect 1702 2000 2322 2016
rect 1702 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1936 1900 2000
rect 1964 1936 1980 2000
rect 2044 1936 2060 2000
rect 2124 1936 2140 2000
rect 2204 1936 2220 2000
rect 2284 1936 2322 2000
rect 1702 0 2322 1936
rect 4702 84592 5322 87000
rect 4702 84528 4740 84592
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84528 5322 84592
rect 4702 84512 5322 84528
rect 4702 84448 4740 84512
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84448 5322 84512
rect 4702 84432 5322 84448
rect 4702 84368 4740 84432
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84368 5322 84432
rect 4702 84352 5322 84368
rect 4702 84288 4740 84352
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84288 5322 84352
rect 4702 74592 5322 84288
rect 4702 74528 4740 74592
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74528 5322 74592
rect 4702 74512 5322 74528
rect 4702 74448 4740 74512
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74448 5322 74512
rect 4702 74432 5322 74448
rect 4702 74368 4740 74432
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74368 5322 74432
rect 4702 74352 5322 74368
rect 4702 74288 4740 74352
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74288 5322 74352
rect 4702 64592 5322 74288
rect 4702 64528 4740 64592
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64528 5322 64592
rect 4702 64512 5322 64528
rect 4702 64448 4740 64512
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64448 5322 64512
rect 4702 64432 5322 64448
rect 4702 64368 4740 64432
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64368 5322 64432
rect 4702 64352 5322 64368
rect 4702 64288 4740 64352
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64288 5322 64352
rect 4702 54592 5322 64288
rect 4702 54528 4740 54592
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54528 5322 54592
rect 4702 54512 5322 54528
rect 4702 54448 4740 54512
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54448 5322 54512
rect 4702 54432 5322 54448
rect 4702 54368 4740 54432
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54368 5322 54432
rect 4702 54352 5322 54368
rect 4702 54288 4740 54352
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54288 5322 54352
rect 4702 44592 5322 54288
rect 4702 44528 4740 44592
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44528 5322 44592
rect 4702 44512 5322 44528
rect 4702 44448 4740 44512
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44448 5322 44512
rect 4702 44432 5322 44448
rect 4702 44368 4740 44432
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44368 5322 44432
rect 4702 44352 5322 44368
rect 4702 44288 4740 44352
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44288 5322 44352
rect 4702 34592 5322 44288
rect 4702 34528 4740 34592
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34528 5322 34592
rect 4702 34512 5322 34528
rect 4702 34448 4740 34512
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34448 5322 34512
rect 4702 34432 5322 34448
rect 4702 34368 4740 34432
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34368 5322 34432
rect 4702 34352 5322 34368
rect 4702 34288 4740 34352
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34288 5322 34352
rect 4702 24592 5322 34288
rect 4702 24528 4740 24592
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24528 5322 24592
rect 4702 24512 5322 24528
rect 4702 24448 4740 24512
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24448 5322 24512
rect 4702 24432 5322 24448
rect 4702 24368 4740 24432
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24368 5322 24432
rect 4702 24352 5322 24368
rect 4702 24288 4740 24352
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24288 5322 24352
rect 4702 14592 5322 24288
rect 4702 14528 4740 14592
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14528 5322 14592
rect 4702 14512 5322 14528
rect 4702 14448 4740 14512
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14448 5322 14512
rect 4702 14432 5322 14448
rect 4702 14368 4740 14432
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14368 5322 14432
rect 4702 14352 5322 14368
rect 4702 14288 4740 14352
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14288 5322 14352
rect 4702 4592 5322 14288
rect 4702 4528 4740 4592
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 5322 4592
rect 4702 4512 5322 4528
rect 4702 4448 4740 4512
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 5322 4512
rect 4702 4432 5322 4448
rect 4702 4368 4740 4432
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 5322 4432
rect 4702 4352 5322 4368
rect 4702 4288 4740 4352
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 5322 4352
rect 4702 0 5322 4288
rect 7702 82240 8322 87000
rect 7702 82176 7740 82240
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82176 8322 82240
rect 7702 82160 8322 82176
rect 7702 82096 7740 82160
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82096 8322 82160
rect 7702 82080 8322 82096
rect 7702 82016 7740 82080
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82016 8322 82080
rect 7702 82000 8322 82016
rect 7702 81936 7740 82000
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81936 8322 82000
rect 7702 72240 8322 81936
rect 7702 72176 7740 72240
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72176 8322 72240
rect 7702 72160 8322 72176
rect 7702 72096 7740 72160
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72096 8322 72160
rect 7702 72080 8322 72096
rect 7702 72016 7740 72080
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72016 8322 72080
rect 7702 72000 8322 72016
rect 7702 71936 7740 72000
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71936 8322 72000
rect 7702 62240 8322 71936
rect 7702 62176 7740 62240
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62176 8322 62240
rect 7702 62160 8322 62176
rect 7702 62096 7740 62160
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62096 8322 62160
rect 7702 62080 8322 62096
rect 7702 62016 7740 62080
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62016 8322 62080
rect 7702 62000 8322 62016
rect 7702 61936 7740 62000
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61936 8322 62000
rect 7702 52240 8322 61936
rect 7702 52176 7740 52240
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52176 8322 52240
rect 7702 52160 8322 52176
rect 7702 52096 7740 52160
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52096 8322 52160
rect 7702 52080 8322 52096
rect 7702 52016 7740 52080
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52016 8322 52080
rect 7702 52000 8322 52016
rect 7702 51936 7740 52000
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51936 8322 52000
rect 7702 42240 8322 51936
rect 7702 42176 7740 42240
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42176 8322 42240
rect 7702 42160 8322 42176
rect 7702 42096 7740 42160
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42096 8322 42160
rect 7702 42080 8322 42096
rect 7702 42016 7740 42080
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42016 8322 42080
rect 7702 42000 8322 42016
rect 7702 41936 7740 42000
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41936 8322 42000
rect 7702 32240 8322 41936
rect 7702 32176 7740 32240
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32176 8322 32240
rect 7702 32160 8322 32176
rect 7702 32096 7740 32160
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32096 8322 32160
rect 7702 32080 8322 32096
rect 7702 32016 7740 32080
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32016 8322 32080
rect 7702 32000 8322 32016
rect 7702 31936 7740 32000
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31936 8322 32000
rect 7702 22240 8322 31936
rect 7702 22176 7740 22240
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22176 8322 22240
rect 7702 22160 8322 22176
rect 7702 22096 7740 22160
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22096 8322 22160
rect 7702 22080 8322 22096
rect 7702 22016 7740 22080
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22016 8322 22080
rect 7702 22000 8322 22016
rect 7702 21936 7740 22000
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21936 8322 22000
rect 7702 12240 8322 21936
rect 7702 12176 7740 12240
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12176 8322 12240
rect 7702 12160 8322 12176
rect 7702 12096 7740 12160
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12096 8322 12160
rect 7702 12080 8322 12096
rect 7702 12016 7740 12080
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12016 8322 12080
rect 7702 12000 8322 12016
rect 7702 11936 7740 12000
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11936 8322 12000
rect 7702 2240 8322 11936
rect 7702 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2176 8322 2240
rect 7702 2160 8322 2176
rect 7702 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2096 8322 2160
rect 7702 2080 8322 2096
rect 7702 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2016 8322 2080
rect 7702 2000 8322 2016
rect 7702 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1936 8322 2000
rect 7702 0 8322 1936
rect 10702 84592 11322 87000
rect 10702 84528 10740 84592
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84528 11322 84592
rect 10702 84512 11322 84528
rect 10702 84448 10740 84512
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84448 11322 84512
rect 10702 84432 11322 84448
rect 10702 84368 10740 84432
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84368 11322 84432
rect 10702 84352 11322 84368
rect 10702 84288 10740 84352
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84288 11322 84352
rect 10702 74592 11322 84288
rect 10702 74528 10740 74592
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74528 11322 74592
rect 10702 74512 11322 74528
rect 10702 74448 10740 74512
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74448 11322 74512
rect 10702 74432 11322 74448
rect 10702 74368 10740 74432
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74368 11322 74432
rect 10702 74352 11322 74368
rect 10702 74288 10740 74352
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74288 11322 74352
rect 10702 64592 11322 74288
rect 10702 64528 10740 64592
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64528 11322 64592
rect 10702 64512 11322 64528
rect 10702 64448 10740 64512
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64448 11322 64512
rect 10702 64432 11322 64448
rect 10702 64368 10740 64432
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64368 11322 64432
rect 10702 64352 11322 64368
rect 10702 64288 10740 64352
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64288 11322 64352
rect 10702 54592 11322 64288
rect 10702 54528 10740 54592
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54528 11322 54592
rect 10702 54512 11322 54528
rect 10702 54448 10740 54512
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54448 11322 54512
rect 10702 54432 11322 54448
rect 10702 54368 10740 54432
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54368 11322 54432
rect 10702 54352 11322 54368
rect 10702 54288 10740 54352
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54288 11322 54352
rect 10702 44592 11322 54288
rect 10702 44528 10740 44592
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44528 11322 44592
rect 10702 44512 11322 44528
rect 10702 44448 10740 44512
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44448 11322 44512
rect 10702 44432 11322 44448
rect 10702 44368 10740 44432
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44368 11322 44432
rect 10702 44352 11322 44368
rect 10702 44288 10740 44352
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44288 11322 44352
rect 10702 34592 11322 44288
rect 10702 34528 10740 34592
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34528 11322 34592
rect 10702 34512 11322 34528
rect 10702 34448 10740 34512
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34448 11322 34512
rect 10702 34432 11322 34448
rect 10702 34368 10740 34432
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34368 11322 34432
rect 10702 34352 11322 34368
rect 10702 34288 10740 34352
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34288 11322 34352
rect 10702 24592 11322 34288
rect 10702 24528 10740 24592
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24528 11322 24592
rect 10702 24512 11322 24528
rect 10702 24448 10740 24512
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24448 11322 24512
rect 10702 24432 11322 24448
rect 10702 24368 10740 24432
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24368 11322 24432
rect 10702 24352 11322 24368
rect 10702 24288 10740 24352
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24288 11322 24352
rect 10702 14592 11322 24288
rect 10702 14528 10740 14592
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14528 11322 14592
rect 10702 14512 11322 14528
rect 10702 14448 10740 14512
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14448 11322 14512
rect 10702 14432 11322 14448
rect 10702 14368 10740 14432
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14368 11322 14432
rect 10702 14352 11322 14368
rect 10702 14288 10740 14352
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14288 11322 14352
rect 10702 4592 11322 14288
rect 10702 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4528 11322 4592
rect 10702 4512 11322 4528
rect 10702 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4448 11322 4512
rect 10702 4432 11322 4448
rect 10702 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4368 11322 4432
rect 10702 4352 11322 4368
rect 10702 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4288 11322 4352
rect 10702 0 11322 4288
rect 13702 82240 14322 87000
rect 13702 82176 13740 82240
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82176 14220 82240
rect 14284 82176 14322 82240
rect 13702 82160 14322 82176
rect 13702 82096 13740 82160
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82096 14220 82160
rect 14284 82096 14322 82160
rect 13702 82080 14322 82096
rect 13702 82016 13740 82080
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82016 14220 82080
rect 14284 82016 14322 82080
rect 13702 82000 14322 82016
rect 13702 81936 13740 82000
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81936 14220 82000
rect 14284 81936 14322 82000
rect 13702 72240 14322 81936
rect 13702 72176 13740 72240
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72176 14220 72240
rect 14284 72176 14322 72240
rect 13702 72160 14322 72176
rect 13702 72096 13740 72160
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72096 14220 72160
rect 14284 72096 14322 72160
rect 13702 72080 14322 72096
rect 13702 72016 13740 72080
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72016 14220 72080
rect 14284 72016 14322 72080
rect 13702 72000 14322 72016
rect 13702 71936 13740 72000
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71936 14220 72000
rect 14284 71936 14322 72000
rect 13702 62240 14322 71936
rect 13702 62176 13740 62240
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62176 14220 62240
rect 14284 62176 14322 62240
rect 13702 62160 14322 62176
rect 13702 62096 13740 62160
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62096 14220 62160
rect 14284 62096 14322 62160
rect 13702 62080 14322 62096
rect 13702 62016 13740 62080
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62016 14220 62080
rect 14284 62016 14322 62080
rect 13702 62000 14322 62016
rect 13702 61936 13740 62000
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61936 14220 62000
rect 14284 61936 14322 62000
rect 13702 52240 14322 61936
rect 13702 52176 13740 52240
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52176 14220 52240
rect 14284 52176 14322 52240
rect 13702 52160 14322 52176
rect 13702 52096 13740 52160
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52096 14220 52160
rect 14284 52096 14322 52160
rect 13702 52080 14322 52096
rect 13702 52016 13740 52080
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52016 14220 52080
rect 14284 52016 14322 52080
rect 13702 52000 14322 52016
rect 13702 51936 13740 52000
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51936 14220 52000
rect 14284 51936 14322 52000
rect 13702 42240 14322 51936
rect 13702 42176 13740 42240
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42176 14220 42240
rect 14284 42176 14322 42240
rect 13702 42160 14322 42176
rect 13702 42096 13740 42160
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42096 14220 42160
rect 14284 42096 14322 42160
rect 13702 42080 14322 42096
rect 13702 42016 13740 42080
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42016 14220 42080
rect 14284 42016 14322 42080
rect 13702 42000 14322 42016
rect 13702 41936 13740 42000
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41936 14220 42000
rect 14284 41936 14322 42000
rect 13702 32240 14322 41936
rect 13702 32176 13740 32240
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32176 14220 32240
rect 14284 32176 14322 32240
rect 13702 32160 14322 32176
rect 13702 32096 13740 32160
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32096 14220 32160
rect 14284 32096 14322 32160
rect 13702 32080 14322 32096
rect 13702 32016 13740 32080
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32016 14220 32080
rect 14284 32016 14322 32080
rect 13702 32000 14322 32016
rect 13702 31936 13740 32000
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31936 14220 32000
rect 14284 31936 14322 32000
rect 13702 22240 14322 31936
rect 13702 22176 13740 22240
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22176 14220 22240
rect 14284 22176 14322 22240
rect 13702 22160 14322 22176
rect 13702 22096 13740 22160
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22096 14220 22160
rect 14284 22096 14322 22160
rect 13702 22080 14322 22096
rect 13702 22016 13740 22080
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22016 14220 22080
rect 14284 22016 14322 22080
rect 13702 22000 14322 22016
rect 13702 21936 13740 22000
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21936 14220 22000
rect 14284 21936 14322 22000
rect 13702 12240 14322 21936
rect 13702 12176 13740 12240
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12176 14220 12240
rect 14284 12176 14322 12240
rect 13702 12160 14322 12176
rect 13702 12096 13740 12160
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12096 14220 12160
rect 14284 12096 14322 12160
rect 13702 12080 14322 12096
rect 13702 12016 13740 12080
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12016 14220 12080
rect 14284 12016 14322 12080
rect 13702 12000 14322 12016
rect 13702 11936 13740 12000
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11936 14220 12000
rect 14284 11936 14322 12000
rect 13702 2240 14322 11936
rect 13702 2176 13740 2240
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 14322 2240
rect 13702 2160 14322 2176
rect 13702 2096 13740 2160
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 14322 2160
rect 13702 2080 14322 2096
rect 13702 2016 13740 2080
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 14322 2080
rect 13702 2000 14322 2016
rect 13702 1936 13740 2000
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 14322 2000
rect 13702 0 14322 1936
rect 16702 84592 17322 87000
rect 16702 84528 16740 84592
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84528 17140 84592
rect 17204 84528 17220 84592
rect 17284 84528 17322 84592
rect 16702 84512 17322 84528
rect 16702 84448 16740 84512
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84448 17140 84512
rect 17204 84448 17220 84512
rect 17284 84448 17322 84512
rect 16702 84432 17322 84448
rect 16702 84368 16740 84432
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84368 17140 84432
rect 17204 84368 17220 84432
rect 17284 84368 17322 84432
rect 16702 84352 17322 84368
rect 16702 84288 16740 84352
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84288 17140 84352
rect 17204 84288 17220 84352
rect 17284 84288 17322 84352
rect 16702 74592 17322 84288
rect 16702 74528 16740 74592
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74528 17140 74592
rect 17204 74528 17220 74592
rect 17284 74528 17322 74592
rect 16702 74512 17322 74528
rect 16702 74448 16740 74512
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74448 17140 74512
rect 17204 74448 17220 74512
rect 17284 74448 17322 74512
rect 16702 74432 17322 74448
rect 16702 74368 16740 74432
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74368 17140 74432
rect 17204 74368 17220 74432
rect 17284 74368 17322 74432
rect 16702 74352 17322 74368
rect 16702 74288 16740 74352
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74288 17140 74352
rect 17204 74288 17220 74352
rect 17284 74288 17322 74352
rect 16702 64592 17322 74288
rect 16702 64528 16740 64592
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64528 17140 64592
rect 17204 64528 17220 64592
rect 17284 64528 17322 64592
rect 16702 64512 17322 64528
rect 16702 64448 16740 64512
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64448 17140 64512
rect 17204 64448 17220 64512
rect 17284 64448 17322 64512
rect 16702 64432 17322 64448
rect 16702 64368 16740 64432
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64368 17140 64432
rect 17204 64368 17220 64432
rect 17284 64368 17322 64432
rect 16702 64352 17322 64368
rect 16702 64288 16740 64352
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64288 17140 64352
rect 17204 64288 17220 64352
rect 17284 64288 17322 64352
rect 16702 54592 17322 64288
rect 16702 54528 16740 54592
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54528 17140 54592
rect 17204 54528 17220 54592
rect 17284 54528 17322 54592
rect 16702 54512 17322 54528
rect 16702 54448 16740 54512
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54448 17140 54512
rect 17204 54448 17220 54512
rect 17284 54448 17322 54512
rect 16702 54432 17322 54448
rect 16702 54368 16740 54432
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54368 17140 54432
rect 17204 54368 17220 54432
rect 17284 54368 17322 54432
rect 16702 54352 17322 54368
rect 16702 54288 16740 54352
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54288 17140 54352
rect 17204 54288 17220 54352
rect 17284 54288 17322 54352
rect 16702 44592 17322 54288
rect 16702 44528 16740 44592
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44528 17140 44592
rect 17204 44528 17220 44592
rect 17284 44528 17322 44592
rect 16702 44512 17322 44528
rect 16702 44448 16740 44512
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44448 17140 44512
rect 17204 44448 17220 44512
rect 17284 44448 17322 44512
rect 16702 44432 17322 44448
rect 16702 44368 16740 44432
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44368 17140 44432
rect 17204 44368 17220 44432
rect 17284 44368 17322 44432
rect 16702 44352 17322 44368
rect 16702 44288 16740 44352
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44288 17140 44352
rect 17204 44288 17220 44352
rect 17284 44288 17322 44352
rect 16702 34592 17322 44288
rect 16702 34528 16740 34592
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34528 17140 34592
rect 17204 34528 17220 34592
rect 17284 34528 17322 34592
rect 16702 34512 17322 34528
rect 16702 34448 16740 34512
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34448 17140 34512
rect 17204 34448 17220 34512
rect 17284 34448 17322 34512
rect 16702 34432 17322 34448
rect 16702 34368 16740 34432
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34368 17140 34432
rect 17204 34368 17220 34432
rect 17284 34368 17322 34432
rect 16702 34352 17322 34368
rect 16702 34288 16740 34352
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34288 17140 34352
rect 17204 34288 17220 34352
rect 17284 34288 17322 34352
rect 16702 24592 17322 34288
rect 16702 24528 16740 24592
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24528 17140 24592
rect 17204 24528 17220 24592
rect 17284 24528 17322 24592
rect 16702 24512 17322 24528
rect 16702 24448 16740 24512
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24448 17140 24512
rect 17204 24448 17220 24512
rect 17284 24448 17322 24512
rect 16702 24432 17322 24448
rect 16702 24368 16740 24432
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24368 17140 24432
rect 17204 24368 17220 24432
rect 17284 24368 17322 24432
rect 16702 24352 17322 24368
rect 16702 24288 16740 24352
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24288 17140 24352
rect 17204 24288 17220 24352
rect 17284 24288 17322 24352
rect 16702 14592 17322 24288
rect 16702 14528 16740 14592
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14528 17140 14592
rect 17204 14528 17220 14592
rect 17284 14528 17322 14592
rect 16702 14512 17322 14528
rect 16702 14448 16740 14512
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14448 17140 14512
rect 17204 14448 17220 14512
rect 17284 14448 17322 14512
rect 16702 14432 17322 14448
rect 16702 14368 16740 14432
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14368 17140 14432
rect 17204 14368 17220 14432
rect 17284 14368 17322 14432
rect 16702 14352 17322 14368
rect 16702 14288 16740 14352
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14288 17140 14352
rect 17204 14288 17220 14352
rect 17284 14288 17322 14352
rect 16702 4592 17322 14288
rect 16702 4528 16740 4592
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 17322 4592
rect 16702 4512 17322 4528
rect 16702 4448 16740 4512
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 17322 4512
rect 16702 4432 17322 4448
rect 16702 4368 16740 4432
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 17322 4432
rect 16702 4352 17322 4368
rect 16702 4288 16740 4352
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 17322 4352
rect 16702 0 17322 4288
rect 19702 82240 20322 87000
rect 19702 82176 19740 82240
rect 19804 82176 19820 82240
rect 19884 82176 19900 82240
rect 19964 82176 19980 82240
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82176 20322 82240
rect 19702 82160 20322 82176
rect 19702 82096 19740 82160
rect 19804 82096 19820 82160
rect 19884 82096 19900 82160
rect 19964 82096 19980 82160
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82096 20322 82160
rect 19702 82080 20322 82096
rect 19702 82016 19740 82080
rect 19804 82016 19820 82080
rect 19884 82016 19900 82080
rect 19964 82016 19980 82080
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82016 20322 82080
rect 19702 82000 20322 82016
rect 19702 81936 19740 82000
rect 19804 81936 19820 82000
rect 19884 81936 19900 82000
rect 19964 81936 19980 82000
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81936 20322 82000
rect 19702 72240 20322 81936
rect 19702 72176 19740 72240
rect 19804 72176 19820 72240
rect 19884 72176 19900 72240
rect 19964 72176 19980 72240
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72176 20322 72240
rect 19702 72160 20322 72176
rect 19702 72096 19740 72160
rect 19804 72096 19820 72160
rect 19884 72096 19900 72160
rect 19964 72096 19980 72160
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72096 20322 72160
rect 19702 72080 20322 72096
rect 19702 72016 19740 72080
rect 19804 72016 19820 72080
rect 19884 72016 19900 72080
rect 19964 72016 19980 72080
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72016 20322 72080
rect 19702 72000 20322 72016
rect 19702 71936 19740 72000
rect 19804 71936 19820 72000
rect 19884 71936 19900 72000
rect 19964 71936 19980 72000
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71936 20322 72000
rect 19702 62240 20322 71936
rect 19702 62176 19740 62240
rect 19804 62176 19820 62240
rect 19884 62176 19900 62240
rect 19964 62176 19980 62240
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62176 20322 62240
rect 19702 62160 20322 62176
rect 19702 62096 19740 62160
rect 19804 62096 19820 62160
rect 19884 62096 19900 62160
rect 19964 62096 19980 62160
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62096 20322 62160
rect 19702 62080 20322 62096
rect 19702 62016 19740 62080
rect 19804 62016 19820 62080
rect 19884 62016 19900 62080
rect 19964 62016 19980 62080
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62016 20322 62080
rect 19702 62000 20322 62016
rect 19702 61936 19740 62000
rect 19804 61936 19820 62000
rect 19884 61936 19900 62000
rect 19964 61936 19980 62000
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61936 20322 62000
rect 19702 52240 20322 61936
rect 19702 52176 19740 52240
rect 19804 52176 19820 52240
rect 19884 52176 19900 52240
rect 19964 52176 19980 52240
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52176 20322 52240
rect 19702 52160 20322 52176
rect 19702 52096 19740 52160
rect 19804 52096 19820 52160
rect 19884 52096 19900 52160
rect 19964 52096 19980 52160
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52096 20322 52160
rect 19702 52080 20322 52096
rect 19702 52016 19740 52080
rect 19804 52016 19820 52080
rect 19884 52016 19900 52080
rect 19964 52016 19980 52080
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52016 20322 52080
rect 19702 52000 20322 52016
rect 19702 51936 19740 52000
rect 19804 51936 19820 52000
rect 19884 51936 19900 52000
rect 19964 51936 19980 52000
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51936 20322 52000
rect 19702 42240 20322 51936
rect 19702 42176 19740 42240
rect 19804 42176 19820 42240
rect 19884 42176 19900 42240
rect 19964 42176 19980 42240
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42176 20322 42240
rect 19702 42160 20322 42176
rect 19702 42096 19740 42160
rect 19804 42096 19820 42160
rect 19884 42096 19900 42160
rect 19964 42096 19980 42160
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42096 20322 42160
rect 19702 42080 20322 42096
rect 19702 42016 19740 42080
rect 19804 42016 19820 42080
rect 19884 42016 19900 42080
rect 19964 42016 19980 42080
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42016 20322 42080
rect 19702 42000 20322 42016
rect 19702 41936 19740 42000
rect 19804 41936 19820 42000
rect 19884 41936 19900 42000
rect 19964 41936 19980 42000
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41936 20322 42000
rect 19702 32240 20322 41936
rect 19702 32176 19740 32240
rect 19804 32176 19820 32240
rect 19884 32176 19900 32240
rect 19964 32176 19980 32240
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32176 20322 32240
rect 19702 32160 20322 32176
rect 19702 32096 19740 32160
rect 19804 32096 19820 32160
rect 19884 32096 19900 32160
rect 19964 32096 19980 32160
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32096 20322 32160
rect 19702 32080 20322 32096
rect 19702 32016 19740 32080
rect 19804 32016 19820 32080
rect 19884 32016 19900 32080
rect 19964 32016 19980 32080
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32016 20322 32080
rect 19702 32000 20322 32016
rect 19702 31936 19740 32000
rect 19804 31936 19820 32000
rect 19884 31936 19900 32000
rect 19964 31936 19980 32000
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31936 20322 32000
rect 19702 22240 20322 31936
rect 19702 22176 19740 22240
rect 19804 22176 19820 22240
rect 19884 22176 19900 22240
rect 19964 22176 19980 22240
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22176 20322 22240
rect 19702 22160 20322 22176
rect 19702 22096 19740 22160
rect 19804 22096 19820 22160
rect 19884 22096 19900 22160
rect 19964 22096 19980 22160
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22096 20322 22160
rect 19702 22080 20322 22096
rect 19702 22016 19740 22080
rect 19804 22016 19820 22080
rect 19884 22016 19900 22080
rect 19964 22016 19980 22080
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22016 20322 22080
rect 19702 22000 20322 22016
rect 19702 21936 19740 22000
rect 19804 21936 19820 22000
rect 19884 21936 19900 22000
rect 19964 21936 19980 22000
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21936 20322 22000
rect 19702 12240 20322 21936
rect 19702 12176 19740 12240
rect 19804 12176 19820 12240
rect 19884 12176 19900 12240
rect 19964 12176 19980 12240
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12176 20322 12240
rect 19702 12160 20322 12176
rect 19702 12096 19740 12160
rect 19804 12096 19820 12160
rect 19884 12096 19900 12160
rect 19964 12096 19980 12160
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12096 20322 12160
rect 19702 12080 20322 12096
rect 19702 12016 19740 12080
rect 19804 12016 19820 12080
rect 19884 12016 19900 12080
rect 19964 12016 19980 12080
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12016 20322 12080
rect 19702 12000 20322 12016
rect 19702 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11936 20322 12000
rect 19702 2240 20322 11936
rect 19702 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2176 20322 2240
rect 19702 2160 20322 2176
rect 19702 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2096 20322 2160
rect 19702 2080 20322 2096
rect 19702 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2016 20322 2080
rect 19702 2000 20322 2016
rect 19702 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1936 20322 2000
rect 19702 0 20322 1936
rect 22702 84592 23322 87000
rect 22702 84528 22740 84592
rect 22804 84528 22820 84592
rect 22884 84528 22900 84592
rect 22964 84528 22980 84592
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84528 23322 84592
rect 22702 84512 23322 84528
rect 22702 84448 22740 84512
rect 22804 84448 22820 84512
rect 22884 84448 22900 84512
rect 22964 84448 22980 84512
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84448 23322 84512
rect 22702 84432 23322 84448
rect 22702 84368 22740 84432
rect 22804 84368 22820 84432
rect 22884 84368 22900 84432
rect 22964 84368 22980 84432
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84368 23322 84432
rect 22702 84352 23322 84368
rect 22702 84288 22740 84352
rect 22804 84288 22820 84352
rect 22884 84288 22900 84352
rect 22964 84288 22980 84352
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84288 23322 84352
rect 22702 74592 23322 84288
rect 22702 74528 22740 74592
rect 22804 74528 22820 74592
rect 22884 74528 22900 74592
rect 22964 74528 22980 74592
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74528 23322 74592
rect 22702 74512 23322 74528
rect 22702 74448 22740 74512
rect 22804 74448 22820 74512
rect 22884 74448 22900 74512
rect 22964 74448 22980 74512
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74448 23322 74512
rect 22702 74432 23322 74448
rect 22702 74368 22740 74432
rect 22804 74368 22820 74432
rect 22884 74368 22900 74432
rect 22964 74368 22980 74432
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74368 23322 74432
rect 22702 74352 23322 74368
rect 22702 74288 22740 74352
rect 22804 74288 22820 74352
rect 22884 74288 22900 74352
rect 22964 74288 22980 74352
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74288 23322 74352
rect 22702 64592 23322 74288
rect 22702 64528 22740 64592
rect 22804 64528 22820 64592
rect 22884 64528 22900 64592
rect 22964 64528 22980 64592
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64528 23322 64592
rect 22702 64512 23322 64528
rect 22702 64448 22740 64512
rect 22804 64448 22820 64512
rect 22884 64448 22900 64512
rect 22964 64448 22980 64512
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64448 23322 64512
rect 22702 64432 23322 64448
rect 22702 64368 22740 64432
rect 22804 64368 22820 64432
rect 22884 64368 22900 64432
rect 22964 64368 22980 64432
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64368 23322 64432
rect 22702 64352 23322 64368
rect 22702 64288 22740 64352
rect 22804 64288 22820 64352
rect 22884 64288 22900 64352
rect 22964 64288 22980 64352
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64288 23322 64352
rect 22702 54592 23322 64288
rect 22702 54528 22740 54592
rect 22804 54528 22820 54592
rect 22884 54528 22900 54592
rect 22964 54528 22980 54592
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54528 23322 54592
rect 22702 54512 23322 54528
rect 22702 54448 22740 54512
rect 22804 54448 22820 54512
rect 22884 54448 22900 54512
rect 22964 54448 22980 54512
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54448 23322 54512
rect 22702 54432 23322 54448
rect 22702 54368 22740 54432
rect 22804 54368 22820 54432
rect 22884 54368 22900 54432
rect 22964 54368 22980 54432
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54368 23322 54432
rect 22702 54352 23322 54368
rect 22702 54288 22740 54352
rect 22804 54288 22820 54352
rect 22884 54288 22900 54352
rect 22964 54288 22980 54352
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54288 23322 54352
rect 22702 44592 23322 54288
rect 22702 44528 22740 44592
rect 22804 44528 22820 44592
rect 22884 44528 22900 44592
rect 22964 44528 22980 44592
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44528 23322 44592
rect 22702 44512 23322 44528
rect 22702 44448 22740 44512
rect 22804 44448 22820 44512
rect 22884 44448 22900 44512
rect 22964 44448 22980 44512
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44448 23322 44512
rect 22702 44432 23322 44448
rect 22702 44368 22740 44432
rect 22804 44368 22820 44432
rect 22884 44368 22900 44432
rect 22964 44368 22980 44432
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44368 23322 44432
rect 22702 44352 23322 44368
rect 22702 44288 22740 44352
rect 22804 44288 22820 44352
rect 22884 44288 22900 44352
rect 22964 44288 22980 44352
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44288 23322 44352
rect 22702 34592 23322 44288
rect 22702 34528 22740 34592
rect 22804 34528 22820 34592
rect 22884 34528 22900 34592
rect 22964 34528 22980 34592
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34528 23322 34592
rect 22702 34512 23322 34528
rect 22702 34448 22740 34512
rect 22804 34448 22820 34512
rect 22884 34448 22900 34512
rect 22964 34448 22980 34512
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34448 23322 34512
rect 22702 34432 23322 34448
rect 22702 34368 22740 34432
rect 22804 34368 22820 34432
rect 22884 34368 22900 34432
rect 22964 34368 22980 34432
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34368 23322 34432
rect 22702 34352 23322 34368
rect 22702 34288 22740 34352
rect 22804 34288 22820 34352
rect 22884 34288 22900 34352
rect 22964 34288 22980 34352
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34288 23322 34352
rect 22702 24592 23322 34288
rect 22702 24528 22740 24592
rect 22804 24528 22820 24592
rect 22884 24528 22900 24592
rect 22964 24528 22980 24592
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24528 23322 24592
rect 22702 24512 23322 24528
rect 22702 24448 22740 24512
rect 22804 24448 22820 24512
rect 22884 24448 22900 24512
rect 22964 24448 22980 24512
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24448 23322 24512
rect 22702 24432 23322 24448
rect 22702 24368 22740 24432
rect 22804 24368 22820 24432
rect 22884 24368 22900 24432
rect 22964 24368 22980 24432
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24368 23322 24432
rect 22702 24352 23322 24368
rect 22702 24288 22740 24352
rect 22804 24288 22820 24352
rect 22884 24288 22900 24352
rect 22964 24288 22980 24352
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24288 23322 24352
rect 22702 14592 23322 24288
rect 22702 14528 22740 14592
rect 22804 14528 22820 14592
rect 22884 14528 22900 14592
rect 22964 14528 22980 14592
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14528 23322 14592
rect 22702 14512 23322 14528
rect 22702 14448 22740 14512
rect 22804 14448 22820 14512
rect 22884 14448 22900 14512
rect 22964 14448 22980 14512
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14448 23322 14512
rect 22702 14432 23322 14448
rect 22702 14368 22740 14432
rect 22804 14368 22820 14432
rect 22884 14368 22900 14432
rect 22964 14368 22980 14432
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14368 23322 14432
rect 22702 14352 23322 14368
rect 22702 14288 22740 14352
rect 22804 14288 22820 14352
rect 22884 14288 22900 14352
rect 22964 14288 22980 14352
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14288 23322 14352
rect 22702 4592 23322 14288
rect 22702 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4528 23322 4592
rect 22702 4512 23322 4528
rect 22702 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4448 23322 4512
rect 22702 4432 23322 4448
rect 22702 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4368 23322 4432
rect 22702 4352 23322 4368
rect 22702 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4288 23322 4352
rect 22702 0 23322 4288
rect 25702 82240 26322 87000
rect 25702 82176 25740 82240
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82176 26322 82240
rect 25702 82160 26322 82176
rect 25702 82096 25740 82160
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82096 26322 82160
rect 25702 82080 26322 82096
rect 25702 82016 25740 82080
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82016 26322 82080
rect 25702 82000 26322 82016
rect 25702 81936 25740 82000
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81936 26322 82000
rect 25702 72240 26322 81936
rect 25702 72176 25740 72240
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72176 26322 72240
rect 25702 72160 26322 72176
rect 25702 72096 25740 72160
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72096 26322 72160
rect 25702 72080 26322 72096
rect 25702 72016 25740 72080
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72016 26322 72080
rect 25702 72000 26322 72016
rect 25702 71936 25740 72000
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71936 26322 72000
rect 25702 62240 26322 71936
rect 25702 62176 25740 62240
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62176 26322 62240
rect 25702 62160 26322 62176
rect 25702 62096 25740 62160
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62096 26322 62160
rect 25702 62080 26322 62096
rect 25702 62016 25740 62080
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62016 26322 62080
rect 25702 62000 26322 62016
rect 25702 61936 25740 62000
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61936 26322 62000
rect 25702 52240 26322 61936
rect 25702 52176 25740 52240
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52176 26322 52240
rect 25702 52160 26322 52176
rect 25702 52096 25740 52160
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52096 26322 52160
rect 25702 52080 26322 52096
rect 25702 52016 25740 52080
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52016 26322 52080
rect 25702 52000 26322 52016
rect 25702 51936 25740 52000
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51936 26322 52000
rect 25702 42240 26322 51936
rect 25702 42176 25740 42240
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42176 26322 42240
rect 25702 42160 26322 42176
rect 25702 42096 25740 42160
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42096 26322 42160
rect 25702 42080 26322 42096
rect 25702 42016 25740 42080
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42016 26322 42080
rect 25702 42000 26322 42016
rect 25702 41936 25740 42000
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41936 26322 42000
rect 25702 32240 26322 41936
rect 25702 32176 25740 32240
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32176 26322 32240
rect 25702 32160 26322 32176
rect 25702 32096 25740 32160
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32096 26322 32160
rect 25702 32080 26322 32096
rect 25702 32016 25740 32080
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32016 26322 32080
rect 25702 32000 26322 32016
rect 25702 31936 25740 32000
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31936 26322 32000
rect 25702 22240 26322 31936
rect 25702 22176 25740 22240
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22176 26322 22240
rect 25702 22160 26322 22176
rect 25702 22096 25740 22160
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22096 26322 22160
rect 25702 22080 26322 22096
rect 25702 22016 25740 22080
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22016 26322 22080
rect 25702 22000 26322 22016
rect 25702 21936 25740 22000
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21936 26322 22000
rect 25702 12240 26322 21936
rect 25702 12176 25740 12240
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12176 26322 12240
rect 25702 12160 26322 12176
rect 25702 12096 25740 12160
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12096 26322 12160
rect 25702 12080 26322 12096
rect 25702 12016 25740 12080
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12016 26322 12080
rect 25702 12000 26322 12016
rect 25702 11936 25740 12000
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11936 26322 12000
rect 25702 2240 26322 11936
rect 25702 2176 25740 2240
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 26322 2240
rect 25702 2160 26322 2176
rect 25702 2096 25740 2160
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 26322 2160
rect 25702 2080 26322 2096
rect 25702 2016 25740 2080
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 26322 2080
rect 25702 2000 26322 2016
rect 25702 1936 25740 2000
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 26322 2000
rect 25702 0 26322 1936
rect 28702 84592 29322 87000
rect 28702 84528 28740 84592
rect 28804 84528 28820 84592
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84528 29322 84592
rect 28702 84512 29322 84528
rect 28702 84448 28740 84512
rect 28804 84448 28820 84512
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84448 29322 84512
rect 28702 84432 29322 84448
rect 28702 84368 28740 84432
rect 28804 84368 28820 84432
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84368 29322 84432
rect 28702 84352 29322 84368
rect 28702 84288 28740 84352
rect 28804 84288 28820 84352
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84288 29322 84352
rect 28702 74592 29322 84288
rect 28702 74528 28740 74592
rect 28804 74528 28820 74592
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74528 29322 74592
rect 28702 74512 29322 74528
rect 28702 74448 28740 74512
rect 28804 74448 28820 74512
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74448 29322 74512
rect 28702 74432 29322 74448
rect 28702 74368 28740 74432
rect 28804 74368 28820 74432
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74368 29322 74432
rect 28702 74352 29322 74368
rect 28702 74288 28740 74352
rect 28804 74288 28820 74352
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74288 29322 74352
rect 28702 64592 29322 74288
rect 28702 64528 28740 64592
rect 28804 64528 28820 64592
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64528 29322 64592
rect 28702 64512 29322 64528
rect 28702 64448 28740 64512
rect 28804 64448 28820 64512
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64448 29322 64512
rect 28702 64432 29322 64448
rect 28702 64368 28740 64432
rect 28804 64368 28820 64432
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64368 29322 64432
rect 28702 64352 29322 64368
rect 28702 64288 28740 64352
rect 28804 64288 28820 64352
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64288 29322 64352
rect 28702 54592 29322 64288
rect 28702 54528 28740 54592
rect 28804 54528 28820 54592
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54528 29322 54592
rect 28702 54512 29322 54528
rect 28702 54448 28740 54512
rect 28804 54448 28820 54512
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54448 29322 54512
rect 28702 54432 29322 54448
rect 28702 54368 28740 54432
rect 28804 54368 28820 54432
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54368 29322 54432
rect 28702 54352 29322 54368
rect 28702 54288 28740 54352
rect 28804 54288 28820 54352
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54288 29322 54352
rect 28702 44592 29322 54288
rect 28702 44528 28740 44592
rect 28804 44528 28820 44592
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44528 29322 44592
rect 28702 44512 29322 44528
rect 28702 44448 28740 44512
rect 28804 44448 28820 44512
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44448 29322 44512
rect 28702 44432 29322 44448
rect 28702 44368 28740 44432
rect 28804 44368 28820 44432
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44368 29322 44432
rect 28702 44352 29322 44368
rect 28702 44288 28740 44352
rect 28804 44288 28820 44352
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44288 29322 44352
rect 28702 34592 29322 44288
rect 28702 34528 28740 34592
rect 28804 34528 28820 34592
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34528 29322 34592
rect 28702 34512 29322 34528
rect 28702 34448 28740 34512
rect 28804 34448 28820 34512
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34448 29322 34512
rect 28702 34432 29322 34448
rect 28702 34368 28740 34432
rect 28804 34368 28820 34432
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34368 29322 34432
rect 28702 34352 29322 34368
rect 28702 34288 28740 34352
rect 28804 34288 28820 34352
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34288 29322 34352
rect 28702 24592 29322 34288
rect 28702 24528 28740 24592
rect 28804 24528 28820 24592
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24528 29322 24592
rect 28702 24512 29322 24528
rect 28702 24448 28740 24512
rect 28804 24448 28820 24512
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24448 29322 24512
rect 28702 24432 29322 24448
rect 28702 24368 28740 24432
rect 28804 24368 28820 24432
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24368 29322 24432
rect 28702 24352 29322 24368
rect 28702 24288 28740 24352
rect 28804 24288 28820 24352
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24288 29322 24352
rect 28702 14592 29322 24288
rect 28702 14528 28740 14592
rect 28804 14528 28820 14592
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14528 29322 14592
rect 28702 14512 29322 14528
rect 28702 14448 28740 14512
rect 28804 14448 28820 14512
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14448 29322 14512
rect 28702 14432 29322 14448
rect 28702 14368 28740 14432
rect 28804 14368 28820 14432
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14368 29322 14432
rect 28702 14352 29322 14368
rect 28702 14288 28740 14352
rect 28804 14288 28820 14352
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14288 29322 14352
rect 28702 4592 29322 14288
rect 28702 4528 28740 4592
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4528 29322 4592
rect 28702 4512 29322 4528
rect 28702 4448 28740 4512
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4448 29322 4512
rect 28702 4432 29322 4448
rect 28702 4368 28740 4432
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4368 29322 4432
rect 28702 4352 29322 4368
rect 28702 4288 28740 4352
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4288 29322 4352
rect 28702 0 29322 4288
rect 31702 82240 32322 87000
rect 31702 82176 31740 82240
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82176 32322 82240
rect 31702 82160 32322 82176
rect 31702 82096 31740 82160
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82096 32322 82160
rect 31702 82080 32322 82096
rect 31702 82016 31740 82080
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82016 32322 82080
rect 31702 82000 32322 82016
rect 31702 81936 31740 82000
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81936 32322 82000
rect 31702 72240 32322 81936
rect 31702 72176 31740 72240
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72176 32322 72240
rect 31702 72160 32322 72176
rect 31702 72096 31740 72160
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72096 32322 72160
rect 31702 72080 32322 72096
rect 31702 72016 31740 72080
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72016 32322 72080
rect 31702 72000 32322 72016
rect 31702 71936 31740 72000
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71936 32322 72000
rect 31702 62240 32322 71936
rect 31702 62176 31740 62240
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62176 32322 62240
rect 31702 62160 32322 62176
rect 31702 62096 31740 62160
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62096 32322 62160
rect 31702 62080 32322 62096
rect 31702 62016 31740 62080
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62016 32322 62080
rect 31702 62000 32322 62016
rect 31702 61936 31740 62000
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61936 32322 62000
rect 31702 52240 32322 61936
rect 31702 52176 31740 52240
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52176 32322 52240
rect 31702 52160 32322 52176
rect 31702 52096 31740 52160
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52096 32322 52160
rect 31702 52080 32322 52096
rect 31702 52016 31740 52080
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52016 32322 52080
rect 31702 52000 32322 52016
rect 31702 51936 31740 52000
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51936 32322 52000
rect 31702 42240 32322 51936
rect 31702 42176 31740 42240
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42176 32322 42240
rect 31702 42160 32322 42176
rect 31702 42096 31740 42160
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42096 32322 42160
rect 31702 42080 32322 42096
rect 31702 42016 31740 42080
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42016 32322 42080
rect 31702 42000 32322 42016
rect 31702 41936 31740 42000
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41936 32322 42000
rect 31702 32240 32322 41936
rect 31702 32176 31740 32240
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32176 32322 32240
rect 31702 32160 32322 32176
rect 31702 32096 31740 32160
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32096 32322 32160
rect 31702 32080 32322 32096
rect 31702 32016 31740 32080
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32016 32322 32080
rect 31702 32000 32322 32016
rect 31702 31936 31740 32000
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31936 32322 32000
rect 31702 22240 32322 31936
rect 31702 22176 31740 22240
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22176 32322 22240
rect 31702 22160 32322 22176
rect 31702 22096 31740 22160
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22096 32322 22160
rect 31702 22080 32322 22096
rect 31702 22016 31740 22080
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22016 32322 22080
rect 31702 22000 32322 22016
rect 31702 21936 31740 22000
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21936 32322 22000
rect 31702 12240 32322 21936
rect 31702 12176 31740 12240
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12176 32322 12240
rect 31702 12160 32322 12176
rect 31702 12096 31740 12160
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12096 32322 12160
rect 31702 12080 32322 12096
rect 31702 12016 31740 12080
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12016 32322 12080
rect 31702 12000 32322 12016
rect 31702 11936 31740 12000
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 32322 12000
rect 31702 2240 32322 11936
rect 31702 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2176 31900 2240
rect 31964 2176 31980 2240
rect 32044 2176 32060 2240
rect 32124 2176 32140 2240
rect 32204 2176 32220 2240
rect 32284 2176 32322 2240
rect 31702 2160 32322 2176
rect 31702 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2096 31900 2160
rect 31964 2096 31980 2160
rect 32044 2096 32060 2160
rect 32124 2096 32140 2160
rect 32204 2096 32220 2160
rect 32284 2096 32322 2160
rect 31702 2080 32322 2096
rect 31702 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2016 31900 2080
rect 31964 2016 31980 2080
rect 32044 2016 32060 2080
rect 32124 2016 32140 2080
rect 32204 2016 32220 2080
rect 32284 2016 32322 2080
rect 31702 2000 32322 2016
rect 31702 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1936 31900 2000
rect 31964 1936 31980 2000
rect 32044 1936 32060 2000
rect 32124 1936 32140 2000
rect 32204 1936 32220 2000
rect 32284 1936 32322 2000
rect 31702 0 32322 1936
rect 34702 84592 35322 87000
rect 34702 84528 34740 84592
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84528 35322 84592
rect 34702 84512 35322 84528
rect 34702 84448 34740 84512
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84448 35322 84512
rect 34702 84432 35322 84448
rect 34702 84368 34740 84432
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84368 35322 84432
rect 34702 84352 35322 84368
rect 34702 84288 34740 84352
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84288 35322 84352
rect 34702 74592 35322 84288
rect 34702 74528 34740 74592
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74528 35322 74592
rect 34702 74512 35322 74528
rect 34702 74448 34740 74512
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74448 35322 74512
rect 34702 74432 35322 74448
rect 34702 74368 34740 74432
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74368 35322 74432
rect 34702 74352 35322 74368
rect 34702 74288 34740 74352
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74288 35322 74352
rect 34702 64592 35322 74288
rect 34702 64528 34740 64592
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64528 35322 64592
rect 34702 64512 35322 64528
rect 34702 64448 34740 64512
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64448 35322 64512
rect 34702 64432 35322 64448
rect 34702 64368 34740 64432
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64368 35322 64432
rect 34702 64352 35322 64368
rect 34702 64288 34740 64352
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64288 35322 64352
rect 34702 54592 35322 64288
rect 34702 54528 34740 54592
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54528 35322 54592
rect 34702 54512 35322 54528
rect 34702 54448 34740 54512
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54448 35322 54512
rect 34702 54432 35322 54448
rect 34702 54368 34740 54432
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54368 35322 54432
rect 34702 54352 35322 54368
rect 34702 54288 34740 54352
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54288 35322 54352
rect 34702 44592 35322 54288
rect 34702 44528 34740 44592
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44528 35322 44592
rect 34702 44512 35322 44528
rect 34702 44448 34740 44512
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44448 35322 44512
rect 34702 44432 35322 44448
rect 34702 44368 34740 44432
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44368 35322 44432
rect 34702 44352 35322 44368
rect 34702 44288 34740 44352
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44288 35322 44352
rect 34702 34592 35322 44288
rect 34702 34528 34740 34592
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34528 35322 34592
rect 34702 34512 35322 34528
rect 34702 34448 34740 34512
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34448 35322 34512
rect 34702 34432 35322 34448
rect 34702 34368 34740 34432
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34368 35322 34432
rect 34702 34352 35322 34368
rect 34702 34288 34740 34352
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34288 35322 34352
rect 34702 24592 35322 34288
rect 34702 24528 34740 24592
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24528 35322 24592
rect 34702 24512 35322 24528
rect 34702 24448 34740 24512
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24448 35322 24512
rect 34702 24432 35322 24448
rect 34702 24368 34740 24432
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24368 35322 24432
rect 34702 24352 35322 24368
rect 34702 24288 34740 24352
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24288 35322 24352
rect 34702 14592 35322 24288
rect 34702 14528 34740 14592
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14528 35322 14592
rect 34702 14512 35322 14528
rect 34702 14448 34740 14512
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14448 35322 14512
rect 34702 14432 35322 14448
rect 34702 14368 34740 14432
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14368 35322 14432
rect 34702 14352 35322 14368
rect 34702 14288 34740 14352
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14288 35322 14352
rect 34702 4592 35322 14288
rect 34702 4528 34740 4592
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 35322 4592
rect 34702 4512 35322 4528
rect 34702 4448 34740 4512
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 35322 4512
rect 34702 4432 35322 4448
rect 34702 4368 34740 4432
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 35322 4432
rect 34702 4352 35322 4368
rect 34702 4288 34740 4352
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 35322 4352
rect 34702 0 35322 4288
rect 37702 82240 38322 87000
rect 37702 82176 37740 82240
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82176 38322 82240
rect 37702 82160 38322 82176
rect 37702 82096 37740 82160
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82096 38322 82160
rect 37702 82080 38322 82096
rect 37702 82016 37740 82080
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82016 38322 82080
rect 37702 82000 38322 82016
rect 37702 81936 37740 82000
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81936 38322 82000
rect 37702 72240 38322 81936
rect 37702 72176 37740 72240
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72176 38322 72240
rect 37702 72160 38322 72176
rect 37702 72096 37740 72160
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72096 38322 72160
rect 37702 72080 38322 72096
rect 37702 72016 37740 72080
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72016 38322 72080
rect 37702 72000 38322 72016
rect 37702 71936 37740 72000
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71936 38322 72000
rect 37702 62240 38322 71936
rect 37702 62176 37740 62240
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62176 38322 62240
rect 37702 62160 38322 62176
rect 37702 62096 37740 62160
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62096 38322 62160
rect 37702 62080 38322 62096
rect 37702 62016 37740 62080
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62016 38322 62080
rect 37702 62000 38322 62016
rect 37702 61936 37740 62000
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61936 38322 62000
rect 37702 52240 38322 61936
rect 37702 52176 37740 52240
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52176 38322 52240
rect 37702 52160 38322 52176
rect 37702 52096 37740 52160
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52096 38322 52160
rect 37702 52080 38322 52096
rect 37702 52016 37740 52080
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52016 38322 52080
rect 37702 52000 38322 52016
rect 37702 51936 37740 52000
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51936 38322 52000
rect 37702 42240 38322 51936
rect 37702 42176 37740 42240
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42176 38322 42240
rect 37702 42160 38322 42176
rect 37702 42096 37740 42160
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42096 38322 42160
rect 37702 42080 38322 42096
rect 37702 42016 37740 42080
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42016 38322 42080
rect 37702 42000 38322 42016
rect 37702 41936 37740 42000
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41936 38322 42000
rect 37702 32240 38322 41936
rect 37702 32176 37740 32240
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32176 38322 32240
rect 37702 32160 38322 32176
rect 37702 32096 37740 32160
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32096 38322 32160
rect 37702 32080 38322 32096
rect 37702 32016 37740 32080
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32016 38322 32080
rect 37702 32000 38322 32016
rect 37702 31936 37740 32000
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31936 38322 32000
rect 37702 22240 38322 31936
rect 37702 22176 37740 22240
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22176 38322 22240
rect 37702 22160 38322 22176
rect 37702 22096 37740 22160
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22096 38322 22160
rect 37702 22080 38322 22096
rect 37702 22016 37740 22080
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22016 38322 22080
rect 37702 22000 38322 22016
rect 37702 21936 37740 22000
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21936 38322 22000
rect 37702 12240 38322 21936
rect 37702 12176 37740 12240
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12176 38322 12240
rect 37702 12160 38322 12176
rect 37702 12096 37740 12160
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12096 38322 12160
rect 37702 12080 38322 12096
rect 37702 12016 37740 12080
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12016 38322 12080
rect 37702 12000 38322 12016
rect 37702 11936 37740 12000
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11936 38322 12000
rect 37702 2240 38322 11936
rect 40702 84592 41322 87000
rect 40702 84528 40740 84592
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84528 41322 84592
rect 40702 84512 41322 84528
rect 40702 84448 40740 84512
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84448 41322 84512
rect 40702 84432 41322 84448
rect 40702 84368 40740 84432
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84368 41322 84432
rect 40702 84352 41322 84368
rect 40702 84288 40740 84352
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84288 41322 84352
rect 40702 74592 41322 84288
rect 40702 74528 40740 74592
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74528 41322 74592
rect 40702 74512 41322 74528
rect 40702 74448 40740 74512
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74448 41322 74512
rect 40702 74432 41322 74448
rect 40702 74368 40740 74432
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74368 41322 74432
rect 40702 74352 41322 74368
rect 40702 74288 40740 74352
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74288 41322 74352
rect 40702 64592 41322 74288
rect 40702 64528 40740 64592
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64528 41322 64592
rect 40702 64512 41322 64528
rect 40702 64448 40740 64512
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64448 41322 64512
rect 40702 64432 41322 64448
rect 40702 64368 40740 64432
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64368 41322 64432
rect 40702 64352 41322 64368
rect 40702 64288 40740 64352
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64288 41322 64352
rect 40702 54592 41322 64288
rect 40702 54528 40740 54592
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54528 41322 54592
rect 40702 54512 41322 54528
rect 40702 54448 40740 54512
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54448 41322 54512
rect 40702 54432 41322 54448
rect 40702 54368 40740 54432
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54368 41322 54432
rect 40702 54352 41322 54368
rect 40702 54288 40740 54352
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54288 41322 54352
rect 40702 44592 41322 54288
rect 40702 44528 40740 44592
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44528 41322 44592
rect 40702 44512 41322 44528
rect 40702 44448 40740 44512
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44448 41322 44512
rect 40702 44432 41322 44448
rect 40702 44368 40740 44432
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44368 41322 44432
rect 40702 44352 41322 44368
rect 40702 44288 40740 44352
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44288 41322 44352
rect 40702 34592 41322 44288
rect 40702 34528 40740 34592
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34528 41322 34592
rect 40702 34512 41322 34528
rect 40702 34448 40740 34512
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34448 41322 34512
rect 40702 34432 41322 34448
rect 40702 34368 40740 34432
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34368 41322 34432
rect 40702 34352 41322 34368
rect 40702 34288 40740 34352
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34288 41322 34352
rect 40702 24592 41322 34288
rect 40702 24528 40740 24592
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24528 41322 24592
rect 40702 24512 41322 24528
rect 40702 24448 40740 24512
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24448 41322 24512
rect 40702 24432 41322 24448
rect 40702 24368 40740 24432
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24368 41322 24432
rect 40702 24352 41322 24368
rect 40702 24288 40740 24352
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24288 41322 24352
rect 40702 14592 41322 24288
rect 40702 14528 40740 14592
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14528 41322 14592
rect 40702 14512 41322 14528
rect 40702 14448 40740 14512
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14448 41322 14512
rect 40702 14432 41322 14448
rect 40702 14368 40740 14432
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14368 41322 14432
rect 40702 14352 41322 14368
rect 40702 14288 40740 14352
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14288 41322 14352
rect 39987 5812 40053 5813
rect 39987 5748 39988 5812
rect 40052 5748 40053 5812
rect 39987 5747 40053 5748
rect 39990 3365 40050 5747
rect 40702 4592 41322 14288
rect 40702 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4528 41322 4592
rect 40702 4512 41322 4528
rect 40702 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4448 41322 4512
rect 40702 4432 41322 4448
rect 40702 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4368 41322 4432
rect 40702 4352 41322 4368
rect 40702 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4288 41322 4352
rect 39987 3364 40053 3365
rect 39987 3300 39988 3364
rect 40052 3300 40053 3364
rect 39987 3299 40053 3300
rect 37702 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2176 38322 2240
rect 37702 2160 38322 2176
rect 37702 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2096 38322 2160
rect 37702 2080 38322 2096
rect 37702 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2016 38322 2080
rect 37702 2000 38322 2016
rect 37702 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1936 38322 2000
rect 37702 0 38322 1936
rect 40702 0 41322 4288
rect 43702 82240 44322 87000
rect 43702 82176 43740 82240
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82176 44322 82240
rect 43702 82160 44322 82176
rect 43702 82096 43740 82160
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82096 44322 82160
rect 43702 82080 44322 82096
rect 43702 82016 43740 82080
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82016 44322 82080
rect 43702 82000 44322 82016
rect 43702 81936 43740 82000
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81936 44322 82000
rect 43702 72240 44322 81936
rect 43702 72176 43740 72240
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72176 44322 72240
rect 43702 72160 44322 72176
rect 43702 72096 43740 72160
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72096 44322 72160
rect 43702 72080 44322 72096
rect 43702 72016 43740 72080
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72016 44322 72080
rect 43702 72000 44322 72016
rect 43702 71936 43740 72000
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71936 44322 72000
rect 43702 62240 44322 71936
rect 43702 62176 43740 62240
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62176 44322 62240
rect 43702 62160 44322 62176
rect 43702 62096 43740 62160
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62096 44322 62160
rect 43702 62080 44322 62096
rect 43702 62016 43740 62080
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62016 44322 62080
rect 43702 62000 44322 62016
rect 43702 61936 43740 62000
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61936 44322 62000
rect 43702 52240 44322 61936
rect 43702 52176 43740 52240
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52176 44322 52240
rect 43702 52160 44322 52176
rect 43702 52096 43740 52160
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52096 44322 52160
rect 43702 52080 44322 52096
rect 43702 52016 43740 52080
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52016 44322 52080
rect 43702 52000 44322 52016
rect 43702 51936 43740 52000
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51936 44322 52000
rect 43702 42240 44322 51936
rect 43702 42176 43740 42240
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42176 44322 42240
rect 43702 42160 44322 42176
rect 43702 42096 43740 42160
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42096 44322 42160
rect 43702 42080 44322 42096
rect 43702 42016 43740 42080
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42016 44322 42080
rect 43702 42000 44322 42016
rect 43702 41936 43740 42000
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41936 44322 42000
rect 43702 32240 44322 41936
rect 43702 32176 43740 32240
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32176 44322 32240
rect 43702 32160 44322 32176
rect 43702 32096 43740 32160
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32096 44322 32160
rect 43702 32080 44322 32096
rect 43702 32016 43740 32080
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32016 44322 32080
rect 43702 32000 44322 32016
rect 43702 31936 43740 32000
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31936 44322 32000
rect 43702 22240 44322 31936
rect 43702 22176 43740 22240
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22176 44322 22240
rect 43702 22160 44322 22176
rect 43702 22096 43740 22160
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22096 44322 22160
rect 43702 22080 44322 22096
rect 43702 22016 43740 22080
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22016 44322 22080
rect 43702 22000 44322 22016
rect 43702 21936 43740 22000
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21936 44322 22000
rect 43702 12240 44322 21936
rect 43702 12176 43740 12240
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12176 44322 12240
rect 43702 12160 44322 12176
rect 43702 12096 43740 12160
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12096 44322 12160
rect 43702 12080 44322 12096
rect 43702 12016 43740 12080
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12016 44322 12080
rect 43702 12000 44322 12016
rect 43702 11936 43740 12000
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11936 44322 12000
rect 43702 2240 44322 11936
rect 43702 2176 43740 2240
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 44322 2240
rect 43702 2160 44322 2176
rect 43702 2096 43740 2160
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 44322 2160
rect 43702 2080 44322 2096
rect 43702 2016 43740 2080
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 44322 2080
rect 43702 2000 44322 2016
rect 43702 1936 43740 2000
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 44322 2000
rect 43702 0 44322 1936
rect 46702 84592 47322 87000
rect 46702 84528 46740 84592
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84528 47322 84592
rect 46702 84512 47322 84528
rect 46702 84448 46740 84512
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84448 47322 84512
rect 46702 84432 47322 84448
rect 46702 84368 46740 84432
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84368 47322 84432
rect 46702 84352 47322 84368
rect 46702 84288 46740 84352
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84288 47322 84352
rect 46702 74592 47322 84288
rect 46702 74528 46740 74592
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74528 47322 74592
rect 46702 74512 47322 74528
rect 46702 74448 46740 74512
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74448 47322 74512
rect 46702 74432 47322 74448
rect 46702 74368 46740 74432
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74368 47322 74432
rect 46702 74352 47322 74368
rect 46702 74288 46740 74352
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74288 47322 74352
rect 46702 64592 47322 74288
rect 46702 64528 46740 64592
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64528 47322 64592
rect 46702 64512 47322 64528
rect 46702 64448 46740 64512
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64448 47322 64512
rect 46702 64432 47322 64448
rect 46702 64368 46740 64432
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64368 47322 64432
rect 46702 64352 47322 64368
rect 46702 64288 46740 64352
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64288 47322 64352
rect 46702 54592 47322 64288
rect 46702 54528 46740 54592
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54528 47322 54592
rect 46702 54512 47322 54528
rect 46702 54448 46740 54512
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54448 47322 54512
rect 46702 54432 47322 54448
rect 46702 54368 46740 54432
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54368 47322 54432
rect 46702 54352 47322 54368
rect 46702 54288 46740 54352
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54288 47322 54352
rect 46702 44592 47322 54288
rect 46702 44528 46740 44592
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44528 47322 44592
rect 46702 44512 47322 44528
rect 46702 44448 46740 44512
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44448 47322 44512
rect 46702 44432 47322 44448
rect 46702 44368 46740 44432
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44368 47322 44432
rect 46702 44352 47322 44368
rect 46702 44288 46740 44352
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44288 47322 44352
rect 46702 34592 47322 44288
rect 46702 34528 46740 34592
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34528 47322 34592
rect 46702 34512 47322 34528
rect 46702 34448 46740 34512
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34448 47322 34512
rect 46702 34432 47322 34448
rect 46702 34368 46740 34432
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34368 47322 34432
rect 46702 34352 47322 34368
rect 46702 34288 46740 34352
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34288 47322 34352
rect 46702 24592 47322 34288
rect 46702 24528 46740 24592
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24528 47322 24592
rect 46702 24512 47322 24528
rect 46702 24448 46740 24512
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24448 47322 24512
rect 46702 24432 47322 24448
rect 46702 24368 46740 24432
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24368 47322 24432
rect 46702 24352 47322 24368
rect 46702 24288 46740 24352
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24288 47322 24352
rect 46702 14592 47322 24288
rect 46702 14528 46740 14592
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14528 47322 14592
rect 46702 14512 47322 14528
rect 46702 14448 46740 14512
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14448 47322 14512
rect 46702 14432 47322 14448
rect 46702 14368 46740 14432
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14368 47322 14432
rect 46702 14352 47322 14368
rect 46702 14288 46740 14352
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14288 47322 14352
rect 46702 4592 47322 14288
rect 46702 4528 46740 4592
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 47322 4592
rect 46702 4512 47322 4528
rect 46702 4448 46740 4512
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 47322 4512
rect 46702 4432 47322 4448
rect 46702 4368 46740 4432
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 47322 4432
rect 46702 4352 47322 4368
rect 46702 4288 46740 4352
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 47322 4352
rect 46702 0 47322 4288
rect 49702 82240 50322 87000
rect 49702 82176 49740 82240
rect 49804 82176 49820 82240
rect 49884 82176 49900 82240
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82176 50322 82240
rect 49702 82160 50322 82176
rect 49702 82096 49740 82160
rect 49804 82096 49820 82160
rect 49884 82096 49900 82160
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82096 50322 82160
rect 49702 82080 50322 82096
rect 49702 82016 49740 82080
rect 49804 82016 49820 82080
rect 49884 82016 49900 82080
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82016 50322 82080
rect 49702 82000 50322 82016
rect 49702 81936 49740 82000
rect 49804 81936 49820 82000
rect 49884 81936 49900 82000
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81936 50322 82000
rect 49702 72240 50322 81936
rect 49702 72176 49740 72240
rect 49804 72176 49820 72240
rect 49884 72176 49900 72240
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72176 50322 72240
rect 49702 72160 50322 72176
rect 49702 72096 49740 72160
rect 49804 72096 49820 72160
rect 49884 72096 49900 72160
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72096 50322 72160
rect 49702 72080 50322 72096
rect 49702 72016 49740 72080
rect 49804 72016 49820 72080
rect 49884 72016 49900 72080
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72016 50322 72080
rect 49702 72000 50322 72016
rect 49702 71936 49740 72000
rect 49804 71936 49820 72000
rect 49884 71936 49900 72000
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71936 50322 72000
rect 49702 62240 50322 71936
rect 49702 62176 49740 62240
rect 49804 62176 49820 62240
rect 49884 62176 49900 62240
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62176 50322 62240
rect 49702 62160 50322 62176
rect 49702 62096 49740 62160
rect 49804 62096 49820 62160
rect 49884 62096 49900 62160
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62096 50322 62160
rect 49702 62080 50322 62096
rect 49702 62016 49740 62080
rect 49804 62016 49820 62080
rect 49884 62016 49900 62080
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62016 50322 62080
rect 49702 62000 50322 62016
rect 49702 61936 49740 62000
rect 49804 61936 49820 62000
rect 49884 61936 49900 62000
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61936 50322 62000
rect 49702 52240 50322 61936
rect 49702 52176 49740 52240
rect 49804 52176 49820 52240
rect 49884 52176 49900 52240
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52176 50322 52240
rect 49702 52160 50322 52176
rect 49702 52096 49740 52160
rect 49804 52096 49820 52160
rect 49884 52096 49900 52160
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52096 50322 52160
rect 49702 52080 50322 52096
rect 49702 52016 49740 52080
rect 49804 52016 49820 52080
rect 49884 52016 49900 52080
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52016 50322 52080
rect 49702 52000 50322 52016
rect 49702 51936 49740 52000
rect 49804 51936 49820 52000
rect 49884 51936 49900 52000
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51936 50322 52000
rect 49702 42240 50322 51936
rect 49702 42176 49740 42240
rect 49804 42176 49820 42240
rect 49884 42176 49900 42240
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42176 50322 42240
rect 49702 42160 50322 42176
rect 49702 42096 49740 42160
rect 49804 42096 49820 42160
rect 49884 42096 49900 42160
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42096 50322 42160
rect 49702 42080 50322 42096
rect 49702 42016 49740 42080
rect 49804 42016 49820 42080
rect 49884 42016 49900 42080
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42016 50322 42080
rect 49702 42000 50322 42016
rect 49702 41936 49740 42000
rect 49804 41936 49820 42000
rect 49884 41936 49900 42000
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41936 50322 42000
rect 49702 32240 50322 41936
rect 49702 32176 49740 32240
rect 49804 32176 49820 32240
rect 49884 32176 49900 32240
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32176 50322 32240
rect 49702 32160 50322 32176
rect 49702 32096 49740 32160
rect 49804 32096 49820 32160
rect 49884 32096 49900 32160
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32096 50322 32160
rect 49702 32080 50322 32096
rect 49702 32016 49740 32080
rect 49804 32016 49820 32080
rect 49884 32016 49900 32080
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32016 50322 32080
rect 49702 32000 50322 32016
rect 49702 31936 49740 32000
rect 49804 31936 49820 32000
rect 49884 31936 49900 32000
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31936 50322 32000
rect 49702 22240 50322 31936
rect 49702 22176 49740 22240
rect 49804 22176 49820 22240
rect 49884 22176 49900 22240
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22176 50322 22240
rect 49702 22160 50322 22176
rect 49702 22096 49740 22160
rect 49804 22096 49820 22160
rect 49884 22096 49900 22160
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22096 50322 22160
rect 49702 22080 50322 22096
rect 49702 22016 49740 22080
rect 49804 22016 49820 22080
rect 49884 22016 49900 22080
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22016 50322 22080
rect 49702 22000 50322 22016
rect 49702 21936 49740 22000
rect 49804 21936 49820 22000
rect 49884 21936 49900 22000
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21936 50322 22000
rect 49702 12240 50322 21936
rect 49702 12176 49740 12240
rect 49804 12176 49820 12240
rect 49884 12176 49900 12240
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12176 50322 12240
rect 49702 12160 50322 12176
rect 49702 12096 49740 12160
rect 49804 12096 49820 12160
rect 49884 12096 49900 12160
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12096 50322 12160
rect 49702 12080 50322 12096
rect 49702 12016 49740 12080
rect 49804 12016 49820 12080
rect 49884 12016 49900 12080
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12016 50322 12080
rect 49702 12000 50322 12016
rect 49702 11936 49740 12000
rect 49804 11936 49820 12000
rect 49884 11936 49900 12000
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11936 50322 12000
rect 49702 2240 50322 11936
rect 49702 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2176 50322 2240
rect 49702 2160 50322 2176
rect 49702 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2096 50322 2160
rect 49702 2080 50322 2096
rect 49702 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2016 50322 2080
rect 49702 2000 50322 2016
rect 49702 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1936 50322 2000
rect 49702 0 50322 1936
rect 52702 84592 53322 87000
rect 52702 84528 52740 84592
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84528 53322 84592
rect 52702 84512 53322 84528
rect 52702 84448 52740 84512
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84448 53322 84512
rect 52702 84432 53322 84448
rect 52702 84368 52740 84432
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84368 53322 84432
rect 52702 84352 53322 84368
rect 52702 84288 52740 84352
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84288 53322 84352
rect 52702 74592 53322 84288
rect 52702 74528 52740 74592
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74528 53322 74592
rect 52702 74512 53322 74528
rect 52702 74448 52740 74512
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74448 53322 74512
rect 52702 74432 53322 74448
rect 52702 74368 52740 74432
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74368 53322 74432
rect 52702 74352 53322 74368
rect 52702 74288 52740 74352
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74288 53322 74352
rect 52702 64592 53322 74288
rect 52702 64528 52740 64592
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64528 53322 64592
rect 52702 64512 53322 64528
rect 52702 64448 52740 64512
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64448 53322 64512
rect 52702 64432 53322 64448
rect 52702 64368 52740 64432
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64368 53322 64432
rect 52702 64352 53322 64368
rect 52702 64288 52740 64352
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64288 53322 64352
rect 52702 54592 53322 64288
rect 52702 54528 52740 54592
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54528 53322 54592
rect 52702 54512 53322 54528
rect 52702 54448 52740 54512
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54448 53322 54512
rect 52702 54432 53322 54448
rect 52702 54368 52740 54432
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54368 53322 54432
rect 52702 54352 53322 54368
rect 52702 54288 52740 54352
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54288 53322 54352
rect 52702 44592 53322 54288
rect 52702 44528 52740 44592
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44528 53322 44592
rect 52702 44512 53322 44528
rect 52702 44448 52740 44512
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44448 53322 44512
rect 52702 44432 53322 44448
rect 52702 44368 52740 44432
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44368 53322 44432
rect 52702 44352 53322 44368
rect 52702 44288 52740 44352
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44288 53322 44352
rect 52702 34592 53322 44288
rect 52702 34528 52740 34592
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34528 53322 34592
rect 52702 34512 53322 34528
rect 52702 34448 52740 34512
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34448 53322 34512
rect 52702 34432 53322 34448
rect 52702 34368 52740 34432
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34368 53322 34432
rect 52702 34352 53322 34368
rect 52702 34288 52740 34352
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34288 53322 34352
rect 52702 24592 53322 34288
rect 52702 24528 52740 24592
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24528 53322 24592
rect 52702 24512 53322 24528
rect 52702 24448 52740 24512
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24448 53322 24512
rect 52702 24432 53322 24448
rect 52702 24368 52740 24432
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24368 53322 24432
rect 52702 24352 53322 24368
rect 52702 24288 52740 24352
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24288 53322 24352
rect 52702 14592 53322 24288
rect 52702 14528 52740 14592
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14528 53322 14592
rect 52702 14512 53322 14528
rect 52702 14448 52740 14512
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14448 53322 14512
rect 52702 14432 53322 14448
rect 52702 14368 52740 14432
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14368 53322 14432
rect 52702 14352 53322 14368
rect 52702 14288 52740 14352
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14288 53322 14352
rect 52702 4592 53322 14288
rect 52702 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4528 53322 4592
rect 52702 4512 53322 4528
rect 52702 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4448 53322 4512
rect 52702 4432 53322 4448
rect 52702 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4368 53322 4432
rect 52702 4352 53322 4368
rect 52702 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4288 53322 4352
rect 52702 0 53322 4288
rect 55702 82240 56322 87000
rect 55702 82176 55740 82240
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82176 56322 82240
rect 55702 82160 56322 82176
rect 55702 82096 55740 82160
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82096 56322 82160
rect 55702 82080 56322 82096
rect 55702 82016 55740 82080
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82016 56322 82080
rect 55702 82000 56322 82016
rect 55702 81936 55740 82000
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81936 56322 82000
rect 55702 72240 56322 81936
rect 55702 72176 55740 72240
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72176 56322 72240
rect 55702 72160 56322 72176
rect 55702 72096 55740 72160
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72096 56322 72160
rect 55702 72080 56322 72096
rect 55702 72016 55740 72080
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72016 56322 72080
rect 55702 72000 56322 72016
rect 55702 71936 55740 72000
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71936 56322 72000
rect 55702 62240 56322 71936
rect 55702 62176 55740 62240
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62176 56322 62240
rect 55702 62160 56322 62176
rect 55702 62096 55740 62160
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62096 56322 62160
rect 55702 62080 56322 62096
rect 55702 62016 55740 62080
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62016 56322 62080
rect 55702 62000 56322 62016
rect 55702 61936 55740 62000
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61936 56322 62000
rect 55702 52240 56322 61936
rect 55702 52176 55740 52240
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52176 56322 52240
rect 55702 52160 56322 52176
rect 55702 52096 55740 52160
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52096 56322 52160
rect 55702 52080 56322 52096
rect 55702 52016 55740 52080
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52016 56322 52080
rect 55702 52000 56322 52016
rect 55702 51936 55740 52000
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51936 56322 52000
rect 55702 42240 56322 51936
rect 55702 42176 55740 42240
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42176 56322 42240
rect 55702 42160 56322 42176
rect 55702 42096 55740 42160
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42096 56322 42160
rect 55702 42080 56322 42096
rect 55702 42016 55740 42080
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42016 56322 42080
rect 55702 42000 56322 42016
rect 55702 41936 55740 42000
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41936 56322 42000
rect 55702 32240 56322 41936
rect 55702 32176 55740 32240
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32176 56322 32240
rect 55702 32160 56322 32176
rect 55702 32096 55740 32160
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32096 56322 32160
rect 55702 32080 56322 32096
rect 55702 32016 55740 32080
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32016 56322 32080
rect 55702 32000 56322 32016
rect 55702 31936 55740 32000
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31936 56322 32000
rect 55702 22240 56322 31936
rect 55702 22176 55740 22240
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22176 56322 22240
rect 55702 22160 56322 22176
rect 55702 22096 55740 22160
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22096 56322 22160
rect 55702 22080 56322 22096
rect 55702 22016 55740 22080
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22016 56322 22080
rect 55702 22000 56322 22016
rect 55702 21936 55740 22000
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21936 56322 22000
rect 55702 12240 56322 21936
rect 55702 12176 55740 12240
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12176 56322 12240
rect 55702 12160 56322 12176
rect 55702 12096 55740 12160
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12096 56322 12160
rect 55702 12080 56322 12096
rect 55702 12016 55740 12080
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12016 56322 12080
rect 55702 12000 56322 12016
rect 55702 11936 55740 12000
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11936 56322 12000
rect 55702 2240 56322 11936
rect 55702 2176 55740 2240
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 56322 2240
rect 55702 2160 56322 2176
rect 55702 2096 55740 2160
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 56322 2160
rect 55702 2080 56322 2096
rect 55702 2016 55740 2080
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 56322 2080
rect 55702 2000 56322 2016
rect 55702 1936 55740 2000
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 56322 2000
rect 55702 0 56322 1936
rect 58702 84592 59322 87000
rect 58702 84528 58740 84592
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84528 59060 84592
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84528 59322 84592
rect 58702 84512 59322 84528
rect 58702 84448 58740 84512
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84448 59060 84512
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84448 59322 84512
rect 58702 84432 59322 84448
rect 58702 84368 58740 84432
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84368 59060 84432
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84368 59322 84432
rect 58702 84352 59322 84368
rect 58702 84288 58740 84352
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84288 59060 84352
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84288 59322 84352
rect 58702 74592 59322 84288
rect 58702 74528 58740 74592
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74528 59060 74592
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74528 59322 74592
rect 58702 74512 59322 74528
rect 58702 74448 58740 74512
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74448 59060 74512
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74448 59322 74512
rect 58702 74432 59322 74448
rect 58702 74368 58740 74432
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74368 59060 74432
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74368 59322 74432
rect 58702 74352 59322 74368
rect 58702 74288 58740 74352
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74288 59060 74352
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74288 59322 74352
rect 58702 64592 59322 74288
rect 58702 64528 58740 64592
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64528 59060 64592
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64528 59322 64592
rect 58702 64512 59322 64528
rect 58702 64448 58740 64512
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64448 59060 64512
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64448 59322 64512
rect 58702 64432 59322 64448
rect 58702 64368 58740 64432
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64368 59060 64432
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64368 59322 64432
rect 58702 64352 59322 64368
rect 58702 64288 58740 64352
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64288 59060 64352
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64288 59322 64352
rect 58702 54592 59322 64288
rect 58702 54528 58740 54592
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54528 59060 54592
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54528 59322 54592
rect 58702 54512 59322 54528
rect 58702 54448 58740 54512
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54448 59060 54512
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54448 59322 54512
rect 58702 54432 59322 54448
rect 58702 54368 58740 54432
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54368 59060 54432
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54368 59322 54432
rect 58702 54352 59322 54368
rect 58702 54288 58740 54352
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54288 59060 54352
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54288 59322 54352
rect 58702 44592 59322 54288
rect 58702 44528 58740 44592
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44528 59060 44592
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44528 59322 44592
rect 58702 44512 59322 44528
rect 58702 44448 58740 44512
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44448 59060 44512
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44448 59322 44512
rect 58702 44432 59322 44448
rect 58702 44368 58740 44432
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44368 59060 44432
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44368 59322 44432
rect 58702 44352 59322 44368
rect 58702 44288 58740 44352
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44288 59060 44352
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44288 59322 44352
rect 58702 34592 59322 44288
rect 58702 34528 58740 34592
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34528 59060 34592
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34528 59322 34592
rect 58702 34512 59322 34528
rect 58702 34448 58740 34512
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34448 59060 34512
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34448 59322 34512
rect 58702 34432 59322 34448
rect 58702 34368 58740 34432
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34368 59060 34432
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34368 59322 34432
rect 58702 34352 59322 34368
rect 58702 34288 58740 34352
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34288 59060 34352
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34288 59322 34352
rect 58702 24592 59322 34288
rect 58702 24528 58740 24592
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24528 59060 24592
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24528 59322 24592
rect 58702 24512 59322 24528
rect 58702 24448 58740 24512
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24448 59060 24512
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24448 59322 24512
rect 58702 24432 59322 24448
rect 58702 24368 58740 24432
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24368 59060 24432
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24368 59322 24432
rect 58702 24352 59322 24368
rect 58702 24288 58740 24352
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24288 59060 24352
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24288 59322 24352
rect 58702 14592 59322 24288
rect 58702 14528 58740 14592
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14528 59060 14592
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14528 59322 14592
rect 58702 14512 59322 14528
rect 58702 14448 58740 14512
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14448 59060 14512
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14448 59322 14512
rect 58702 14432 59322 14448
rect 58702 14368 58740 14432
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14368 59060 14432
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14368 59322 14432
rect 58702 14352 59322 14368
rect 58702 14288 58740 14352
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14288 59060 14352
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14288 59322 14352
rect 58702 4592 59322 14288
rect 58702 4528 58740 4592
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4528 59322 4592
rect 58702 4512 59322 4528
rect 58702 4448 58740 4512
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4448 59322 4512
rect 58702 4432 59322 4448
rect 58702 4368 58740 4432
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4368 59322 4432
rect 58702 4352 59322 4368
rect 58702 4288 58740 4352
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4288 59322 4352
rect 58702 0 59322 4288
rect 61702 82240 62322 87000
rect 61702 82176 61740 82240
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82176 62322 82240
rect 61702 82160 62322 82176
rect 61702 82096 61740 82160
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82096 62322 82160
rect 61702 82080 62322 82096
rect 61702 82016 61740 82080
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82016 62322 82080
rect 61702 82000 62322 82016
rect 61702 81936 61740 82000
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81936 62322 82000
rect 61702 72240 62322 81936
rect 61702 72176 61740 72240
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72176 62322 72240
rect 61702 72160 62322 72176
rect 61702 72096 61740 72160
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72096 62322 72160
rect 61702 72080 62322 72096
rect 61702 72016 61740 72080
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72016 62322 72080
rect 61702 72000 62322 72016
rect 61702 71936 61740 72000
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71936 62322 72000
rect 61702 62240 62322 71936
rect 61702 62176 61740 62240
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62176 62322 62240
rect 61702 62160 62322 62176
rect 61702 62096 61740 62160
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62096 62322 62160
rect 61702 62080 62322 62096
rect 61702 62016 61740 62080
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62016 62322 62080
rect 61702 62000 62322 62016
rect 61702 61936 61740 62000
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61936 62322 62000
rect 61702 52240 62322 61936
rect 64702 84592 65322 87000
rect 64702 84528 64740 84592
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 65322 84592
rect 64702 84512 65322 84528
rect 64702 84448 64740 84512
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 65322 84512
rect 64702 84432 65322 84448
rect 64702 84368 64740 84432
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 65322 84432
rect 64702 84352 65322 84368
rect 64702 84288 64740 84352
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 65322 84352
rect 64702 74592 65322 84288
rect 64702 74528 64740 74592
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 65322 74592
rect 64702 74512 65322 74528
rect 64702 74448 64740 74512
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 65322 74512
rect 64702 74432 65322 74448
rect 64702 74368 64740 74432
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 65322 74432
rect 64702 74352 65322 74368
rect 64702 74288 64740 74352
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 65322 74352
rect 64702 64592 65322 74288
rect 64702 64528 64740 64592
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 65322 64592
rect 64702 64512 65322 64528
rect 64702 64448 64740 64512
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 65322 64512
rect 64702 64432 65322 64448
rect 64702 64368 64740 64432
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 65322 64432
rect 64702 64352 65322 64368
rect 64702 64288 64740 64352
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 65322 64352
rect 64702 54592 65322 64288
rect 64702 54528 64740 54592
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 65322 54592
rect 64702 54512 65322 54528
rect 64702 54448 64740 54512
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 65322 54512
rect 64702 54432 65322 54448
rect 64702 54368 64740 54432
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 65322 54432
rect 64702 54352 65322 54368
rect 64702 54288 64740 54352
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 65322 54352
rect 64091 52596 64157 52597
rect 64091 52532 64092 52596
rect 64156 52532 64157 52596
rect 64091 52531 64157 52532
rect 61702 52176 61740 52240
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52176 62322 52240
rect 61702 52160 62322 52176
rect 61702 52096 61740 52160
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52096 62322 52160
rect 61702 52080 62322 52096
rect 61702 52016 61740 52080
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52016 62322 52080
rect 61702 52000 62322 52016
rect 61702 51936 61740 52000
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51936 62322 52000
rect 61702 42240 62322 51936
rect 62987 48788 63053 48789
rect 62987 48724 62988 48788
rect 63052 48724 63053 48788
rect 62987 48723 63053 48724
rect 61702 42176 61740 42240
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42176 62322 42240
rect 61702 42160 62322 42176
rect 61702 42096 61740 42160
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42096 62322 42160
rect 61702 42080 62322 42096
rect 61702 42016 61740 42080
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42016 62322 42080
rect 61702 42000 62322 42016
rect 61702 41936 61740 42000
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41936 62322 42000
rect 61702 32240 62322 41936
rect 61702 32176 61740 32240
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32176 62322 32240
rect 61702 32160 62322 32176
rect 61702 32096 61740 32160
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32096 62322 32160
rect 61702 32080 62322 32096
rect 61702 32016 61740 32080
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32016 62322 32080
rect 61702 32000 62322 32016
rect 61702 31936 61740 32000
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31936 62322 32000
rect 61702 22240 62322 31936
rect 61702 22176 61740 22240
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22176 62322 22240
rect 61702 22160 62322 22176
rect 61702 22096 61740 22160
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22096 62322 22160
rect 61702 22080 62322 22096
rect 61702 22016 61740 22080
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22016 62322 22080
rect 61702 22000 62322 22016
rect 61702 21936 61740 22000
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21936 62322 22000
rect 61702 12240 62322 21936
rect 61702 12176 61740 12240
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12176 62322 12240
rect 61702 12160 62322 12176
rect 61702 12096 61740 12160
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12096 62322 12160
rect 61702 12080 62322 12096
rect 61702 12016 61740 12080
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12016 62322 12080
rect 61702 12000 62322 12016
rect 61702 11936 61740 12000
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11936 62322 12000
rect 61702 2240 62322 11936
rect 62990 7581 63050 48723
rect 63907 47700 63973 47701
rect 63907 47636 63908 47700
rect 63972 47636 63973 47700
rect 63907 47635 63973 47636
rect 63171 26212 63237 26213
rect 63171 26148 63172 26212
rect 63236 26148 63237 26212
rect 63171 26147 63237 26148
rect 62987 7580 63053 7581
rect 62987 7516 62988 7580
rect 63052 7516 63053 7580
rect 62987 7515 63053 7516
rect 63174 5813 63234 26147
rect 63910 19350 63970 47635
rect 63358 19290 63970 19350
rect 63358 11661 63418 19290
rect 63539 16556 63605 16557
rect 63539 16492 63540 16556
rect 63604 16492 63605 16556
rect 63539 16491 63605 16492
rect 63542 11797 63602 16491
rect 63723 14788 63789 14789
rect 63723 14724 63724 14788
rect 63788 14724 63789 14788
rect 63723 14723 63789 14724
rect 63539 11796 63605 11797
rect 63539 11732 63540 11796
rect 63604 11732 63605 11796
rect 63539 11731 63605 11732
rect 63355 11660 63421 11661
rect 63355 11596 63356 11660
rect 63420 11596 63421 11660
rect 63355 11595 63421 11596
rect 63355 10708 63421 10709
rect 63355 10644 63356 10708
rect 63420 10644 63421 10708
rect 63355 10643 63421 10644
rect 63358 7309 63418 10643
rect 63355 7308 63421 7309
rect 63355 7244 63356 7308
rect 63420 7244 63421 7308
rect 63355 7243 63421 7244
rect 63171 5812 63237 5813
rect 63171 5748 63172 5812
rect 63236 5748 63237 5812
rect 63171 5747 63237 5748
rect 63726 4045 63786 14723
rect 64094 12613 64154 52531
rect 64275 50284 64341 50285
rect 64275 50220 64276 50284
rect 64340 50220 64341 50284
rect 64275 50219 64341 50220
rect 64091 12612 64157 12613
rect 64091 12548 64092 12612
rect 64156 12548 64157 12612
rect 64278 12610 64338 50219
rect 64459 48108 64525 48109
rect 64459 48044 64460 48108
rect 64524 48044 64525 48108
rect 64459 48043 64525 48044
rect 64462 14789 64522 48043
rect 64702 44592 65322 54288
rect 64702 44528 64740 44592
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 65322 44592
rect 64702 44512 65322 44528
rect 64702 44448 64740 44512
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 65322 44512
rect 64702 44432 65322 44448
rect 64702 44368 64740 44432
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 65322 44432
rect 64702 44352 65322 44368
rect 64702 44288 64740 44352
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 65322 44352
rect 64702 34592 65322 44288
rect 67702 82240 68322 87000
rect 67702 82176 67740 82240
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82176 68322 82240
rect 67702 82160 68322 82176
rect 67702 82096 67740 82160
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82096 68322 82160
rect 67702 82080 68322 82096
rect 67702 82016 67740 82080
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82016 68322 82080
rect 67702 82000 68322 82016
rect 67702 81936 67740 82000
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81936 68322 82000
rect 67702 72240 68322 81936
rect 67702 72176 67740 72240
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72176 68322 72240
rect 67702 72160 68322 72176
rect 67702 72096 67740 72160
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72096 68322 72160
rect 67702 72080 68322 72096
rect 67702 72016 67740 72080
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72016 68322 72080
rect 67702 72000 68322 72016
rect 67702 71936 67740 72000
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71936 68322 72000
rect 67702 62240 68322 71936
rect 67702 62176 67740 62240
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62176 68322 62240
rect 67702 62160 68322 62176
rect 67702 62096 67740 62160
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62096 68322 62160
rect 67702 62080 68322 62096
rect 67702 62016 67740 62080
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62016 68322 62080
rect 67702 62000 68322 62016
rect 67702 61936 67740 62000
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61936 68322 62000
rect 67702 52240 68322 61936
rect 67702 52176 67740 52240
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52176 68322 52240
rect 67702 52160 68322 52176
rect 67702 52096 67740 52160
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52096 68322 52160
rect 67702 52080 68322 52096
rect 67702 52016 67740 52080
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52016 68322 52080
rect 67702 52000 68322 52016
rect 67702 51936 67740 52000
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51936 68322 52000
rect 67702 42240 68322 51936
rect 67702 42176 67740 42240
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42176 68322 42240
rect 67702 42160 68322 42176
rect 67702 42096 67740 42160
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42096 68322 42160
rect 67702 42080 68322 42096
rect 67702 42016 67740 42080
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42016 68322 42080
rect 67702 42000 68322 42016
rect 67702 41936 67740 42000
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41936 68322 42000
rect 65563 40900 65629 40901
rect 65563 40836 65564 40900
rect 65628 40836 65629 40900
rect 65563 40835 65629 40836
rect 64702 34528 64740 34592
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 65322 34592
rect 64702 34512 65322 34528
rect 64702 34448 64740 34512
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 65322 34512
rect 64702 34432 65322 34448
rect 64702 34368 64740 34432
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 65322 34432
rect 64702 34352 65322 34368
rect 64702 34288 64740 34352
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 65322 34352
rect 64702 24592 65322 34288
rect 64702 24528 64740 24592
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 65322 24592
rect 64702 24512 65322 24528
rect 64702 24448 64740 24512
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 65322 24512
rect 64702 24432 65322 24448
rect 64702 24368 64740 24432
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 65322 24432
rect 64702 24352 65322 24368
rect 64702 24288 64740 24352
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 65322 24352
rect 64459 14788 64525 14789
rect 64459 14724 64460 14788
rect 64524 14724 64525 14788
rect 64459 14723 64525 14724
rect 64702 14592 65322 24288
rect 64702 14528 64740 14592
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 65322 14592
rect 64702 14512 65322 14528
rect 64702 14448 64740 14512
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 65322 14512
rect 64702 14432 65322 14448
rect 64702 14368 64740 14432
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 65322 14432
rect 64702 14352 65322 14368
rect 64702 14288 64740 14352
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 65322 14352
rect 64278 12550 64522 12610
rect 64091 12547 64157 12548
rect 64275 11796 64341 11797
rect 64275 11732 64276 11796
rect 64340 11732 64341 11796
rect 64275 11731 64341 11732
rect 63907 11660 63973 11661
rect 63907 11596 63908 11660
rect 63972 11596 63973 11660
rect 63907 11595 63973 11596
rect 63910 7717 63970 11595
rect 64091 11116 64157 11117
rect 64091 11052 64092 11116
rect 64156 11052 64157 11116
rect 64091 11051 64157 11052
rect 63907 7716 63973 7717
rect 63907 7652 63908 7716
rect 63972 7652 63973 7716
rect 63907 7651 63973 7652
rect 64094 7037 64154 11051
rect 64091 7036 64157 7037
rect 64091 6972 64092 7036
rect 64156 6972 64157 7036
rect 64091 6971 64157 6972
rect 64278 5133 64338 11731
rect 64275 5132 64341 5133
rect 64275 5068 64276 5132
rect 64340 5068 64341 5132
rect 64275 5067 64341 5068
rect 64462 4997 64522 12550
rect 64459 4996 64525 4997
rect 64459 4932 64460 4996
rect 64524 4932 64525 4996
rect 64459 4931 64525 4932
rect 64702 4592 65322 14288
rect 65566 6765 65626 40835
rect 65747 38860 65813 38861
rect 65747 38796 65748 38860
rect 65812 38796 65813 38860
rect 65747 38795 65813 38796
rect 65563 6764 65629 6765
rect 65563 6700 65564 6764
rect 65628 6700 65629 6764
rect 65563 6699 65629 6700
rect 65750 6629 65810 38795
rect 65931 34780 65997 34781
rect 65931 34716 65932 34780
rect 65996 34716 65997 34780
rect 65931 34715 65997 34716
rect 65747 6628 65813 6629
rect 65747 6564 65748 6628
rect 65812 6564 65813 6628
rect 65747 6563 65813 6564
rect 65934 6085 65994 34715
rect 67702 32240 68322 41936
rect 70702 84592 71322 87000
rect 70702 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84528 71322 84592
rect 70702 84512 71322 84528
rect 70702 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84448 71322 84512
rect 70702 84432 71322 84448
rect 70702 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84368 71322 84432
rect 70702 84352 71322 84368
rect 70702 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84288 71322 84352
rect 70702 74592 71322 84288
rect 70702 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74528 71322 74592
rect 70702 74512 71322 74528
rect 70702 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74448 71322 74512
rect 70702 74432 71322 74448
rect 70702 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74368 71322 74432
rect 70702 74352 71322 74368
rect 70702 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74288 71322 74352
rect 70702 64592 71322 74288
rect 70702 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64528 71322 64592
rect 70702 64512 71322 64528
rect 70702 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64448 71322 64512
rect 70702 64432 71322 64448
rect 70702 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64368 71322 64432
rect 70702 64352 71322 64368
rect 70702 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64288 71322 64352
rect 70702 54592 71322 64288
rect 70702 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54528 71322 54592
rect 70702 54512 71322 54528
rect 70702 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54448 71322 54512
rect 70702 54432 71322 54448
rect 70702 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54368 71322 54432
rect 70702 54352 71322 54368
rect 70702 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54288 71322 54352
rect 70702 44592 71322 54288
rect 70702 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44528 71322 44592
rect 70702 44512 71322 44528
rect 70702 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44448 71322 44512
rect 70702 44432 71322 44448
rect 70702 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44368 71322 44432
rect 70702 44352 71322 44368
rect 70702 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44288 71322 44352
rect 70702 34592 71322 44288
rect 70702 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34528 71322 34592
rect 70702 34512 71322 34528
rect 70702 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34448 71322 34512
rect 70702 34432 71322 34448
rect 70702 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34368 71322 34432
rect 70702 34352 71322 34368
rect 70702 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34288 71322 34352
rect 68507 33284 68573 33285
rect 68507 33220 68508 33284
rect 68572 33220 68573 33284
rect 68507 33219 68573 33220
rect 67702 32176 67740 32240
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32176 68322 32240
rect 67702 32160 68322 32176
rect 67702 32096 67740 32160
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32096 68322 32160
rect 67702 32080 68322 32096
rect 67702 32016 67740 32080
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32016 68322 32080
rect 67702 32000 68322 32016
rect 67702 31936 67740 32000
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31936 68322 32000
rect 67403 26484 67469 26485
rect 67403 26420 67404 26484
rect 67468 26420 67469 26484
rect 67403 26419 67469 26420
rect 67406 26077 67466 26419
rect 67403 26076 67469 26077
rect 67403 26012 67404 26076
rect 67468 26012 67469 26076
rect 67403 26011 67469 26012
rect 66483 23628 66549 23629
rect 66483 23564 66484 23628
rect 66548 23564 66549 23628
rect 66483 23563 66549 23564
rect 66299 23492 66365 23493
rect 66299 23428 66300 23492
rect 66364 23428 66365 23492
rect 66299 23427 66365 23428
rect 65931 6084 65997 6085
rect 65931 6020 65932 6084
rect 65996 6020 65997 6084
rect 65931 6019 65997 6020
rect 64702 4528 64740 4592
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 65322 4592
rect 64702 4512 65322 4528
rect 64702 4448 64740 4512
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 65322 4512
rect 64702 4432 65322 4448
rect 64702 4368 64740 4432
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 65322 4432
rect 64702 4352 65322 4368
rect 64702 4288 64740 4352
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 65322 4352
rect 63723 4044 63789 4045
rect 63723 3980 63724 4044
rect 63788 3980 63789 4044
rect 63723 3979 63789 3980
rect 61702 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2176 61900 2240
rect 61964 2176 61980 2240
rect 62044 2176 62060 2240
rect 62124 2176 62140 2240
rect 62204 2176 62220 2240
rect 62284 2176 62322 2240
rect 61702 2160 62322 2176
rect 61702 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2096 61900 2160
rect 61964 2096 61980 2160
rect 62044 2096 62060 2160
rect 62124 2096 62140 2160
rect 62204 2096 62220 2160
rect 62284 2096 62322 2160
rect 61702 2080 62322 2096
rect 61702 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2016 61900 2080
rect 61964 2016 61980 2080
rect 62044 2016 62060 2080
rect 62124 2016 62140 2080
rect 62204 2016 62220 2080
rect 62284 2016 62322 2080
rect 61702 2000 62322 2016
rect 61702 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1936 61900 2000
rect 61964 1936 61980 2000
rect 62044 1936 62060 2000
rect 62124 1936 62140 2000
rect 62204 1936 62220 2000
rect 62284 1936 62322 2000
rect 61702 0 62322 1936
rect 64702 0 65322 4288
rect 66302 3365 66362 23427
rect 66486 6357 66546 23563
rect 66667 22404 66733 22405
rect 66667 22340 66668 22404
rect 66732 22340 66733 22404
rect 66667 22339 66733 22340
rect 66483 6356 66549 6357
rect 66483 6292 66484 6356
rect 66548 6292 66549 6356
rect 66483 6291 66549 6292
rect 66670 4861 66730 22339
rect 67702 22240 68322 31936
rect 67702 22176 67740 22240
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22176 68322 22240
rect 67702 22160 68322 22176
rect 67702 22096 67740 22160
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22096 68322 22160
rect 67702 22080 68322 22096
rect 67702 22016 67740 22080
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22016 68322 22080
rect 67702 22000 68322 22016
rect 67702 21936 67740 22000
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21936 68322 22000
rect 66851 12748 66917 12749
rect 66851 12684 66852 12748
rect 66916 12684 66917 12748
rect 66851 12683 66917 12684
rect 66854 6221 66914 12683
rect 67702 12240 68322 21936
rect 67702 12176 67740 12240
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12176 68322 12240
rect 67702 12160 68322 12176
rect 67702 12096 67740 12160
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12096 68322 12160
rect 67702 12080 68322 12096
rect 67702 12016 67740 12080
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12016 68322 12080
rect 67702 12000 68322 12016
rect 67702 11936 67740 12000
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11936 68322 12000
rect 66851 6220 66917 6221
rect 66851 6156 66852 6220
rect 66916 6156 66917 6220
rect 66851 6155 66917 6156
rect 66667 4860 66733 4861
rect 66667 4796 66668 4860
rect 66732 4796 66733 4860
rect 66667 4795 66733 4796
rect 66299 3364 66365 3365
rect 66299 3300 66300 3364
rect 66364 3300 66365 3364
rect 66299 3299 66365 3300
rect 67702 2240 68322 11936
rect 68510 5677 68570 33219
rect 70702 24592 71322 34288
rect 70702 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24528 71322 24592
rect 70702 24512 71322 24528
rect 70702 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24448 71322 24512
rect 70702 24432 71322 24448
rect 70702 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24368 71322 24432
rect 70702 24352 71322 24368
rect 70702 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24288 71322 24352
rect 70702 14592 71322 24288
rect 70702 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14528 71322 14592
rect 70702 14512 71322 14528
rect 70702 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14448 71322 14512
rect 70702 14432 71322 14448
rect 70702 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14368 71322 14432
rect 70702 14352 71322 14368
rect 70702 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14288 71322 14352
rect 68507 5676 68573 5677
rect 68507 5612 68508 5676
rect 68572 5612 68573 5676
rect 68507 5611 68573 5612
rect 67702 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2176 68322 2240
rect 67702 2160 68322 2176
rect 67702 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2096 68322 2160
rect 67702 2080 68322 2096
rect 67702 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2016 68322 2080
rect 67702 2000 68322 2016
rect 67702 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1936 68322 2000
rect 67702 0 68322 1936
rect 70702 4592 71322 14288
rect 70702 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4528 71322 4592
rect 70702 4512 71322 4528
rect 70702 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4448 71322 4512
rect 70702 4432 71322 4448
rect 70702 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4368 71322 4432
rect 70702 4352 71322 4368
rect 70702 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4288 71322 4352
rect 70702 0 71322 4288
rect 73702 82240 74322 87000
rect 73702 82176 73740 82240
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 74322 82240
rect 73702 82160 74322 82176
rect 73702 82096 73740 82160
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 74322 82160
rect 73702 82080 74322 82096
rect 73702 82016 73740 82080
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 74322 82080
rect 73702 82000 74322 82016
rect 73702 81936 73740 82000
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 74322 82000
rect 73702 72240 74322 81936
rect 73702 72176 73740 72240
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 74322 72240
rect 73702 72160 74322 72176
rect 73702 72096 73740 72160
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 74322 72160
rect 73702 72080 74322 72096
rect 73702 72016 73740 72080
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 74322 72080
rect 73702 72000 74322 72016
rect 73702 71936 73740 72000
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 74322 72000
rect 73702 62240 74322 71936
rect 73702 62176 73740 62240
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 74322 62240
rect 73702 62160 74322 62176
rect 73702 62096 73740 62160
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 74322 62160
rect 73702 62080 74322 62096
rect 73702 62016 73740 62080
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 74322 62080
rect 73702 62000 74322 62016
rect 73702 61936 73740 62000
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 74322 62000
rect 73702 52240 74322 61936
rect 73702 52176 73740 52240
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 74322 52240
rect 73702 52160 74322 52176
rect 73702 52096 73740 52160
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 74322 52160
rect 73702 52080 74322 52096
rect 73702 52016 73740 52080
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 74322 52080
rect 73702 52000 74322 52016
rect 73702 51936 73740 52000
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 74322 52000
rect 73702 42240 74322 51936
rect 73702 42176 73740 42240
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 74322 42240
rect 73702 42160 74322 42176
rect 73702 42096 73740 42160
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 74322 42160
rect 73702 42080 74322 42096
rect 73702 42016 73740 42080
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 74322 42080
rect 73702 42000 74322 42016
rect 73702 41936 73740 42000
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 74322 42000
rect 73702 32240 74322 41936
rect 73702 32176 73740 32240
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 74322 32240
rect 73702 32160 74322 32176
rect 73702 32096 73740 32160
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 74322 32160
rect 73702 32080 74322 32096
rect 73702 32016 73740 32080
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 74322 32080
rect 73702 32000 74322 32016
rect 73702 31936 73740 32000
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 74322 32000
rect 73702 22240 74322 31936
rect 73702 22176 73740 22240
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 74322 22240
rect 73702 22160 74322 22176
rect 73702 22096 73740 22160
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 74322 22160
rect 73702 22080 74322 22096
rect 73702 22016 73740 22080
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 74322 22080
rect 73702 22000 74322 22016
rect 73702 21936 73740 22000
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 74322 22000
rect 73702 12240 74322 21936
rect 73702 12176 73740 12240
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 74322 12240
rect 73702 12160 74322 12176
rect 73702 12096 73740 12160
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 74322 12160
rect 73702 12080 74322 12096
rect 73702 12016 73740 12080
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 74322 12080
rect 73702 12000 74322 12016
rect 73702 11936 73740 12000
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 74322 12000
rect 73702 2240 74322 11936
rect 73702 2176 73740 2240
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 74322 2240
rect 73702 2160 74322 2176
rect 73702 2096 73740 2160
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 74322 2160
rect 73702 2080 74322 2096
rect 73702 2016 73740 2080
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 74322 2080
rect 73702 2000 74322 2016
rect 73702 1936 73740 2000
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 74322 2000
rect 73702 0 74322 1936
use sky130_fd_sc_hd__nor2b_4  _049_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 44436 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _050_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _051_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 30912 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25944 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _053_
timestamp 1704896540
transform -1 0 30360 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1704896540
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _055_
timestamp 1704896540
transform -1 0 29808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp 1704896540
transform -1 0 26772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _057_
timestamp 1704896540
transform -1 0 29164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp 1704896540
transform -1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _059_
timestamp 1704896540
transform -1 0 28520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp 1704896540
transform -1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _061_
timestamp 1704896540
transform 1 0 27048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp 1704896540
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _063_
timestamp 1704896540
transform 1 0 26312 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp 1704896540
transform 1 0 29440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _065_
timestamp 1704896540
transform 1 0 25852 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp 1704896540
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _067_
timestamp 1704896540
transform 1 0 24196 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp 1704896540
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _069_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 35052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _070_
timestamp 1704896540
transform 1 0 25392 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp 1704896540
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _072_
timestamp 1704896540
transform 1 0 24748 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _073_
timestamp 1704896540
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _074_
timestamp 1704896540
transform 1 0 24288 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp 1704896540
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _076_
timestamp 1704896540
transform 1 0 23276 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp 1704896540
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _078_
timestamp 1704896540
transform 1 0 23736 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp 1704896540
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _080_
timestamp 1704896540
transform 1 0 25760 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp 1704896540
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _082_
timestamp 1704896540
transform 1 0 27508 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp 1704896540
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _084_
timestamp 1704896540
transform 1 0 44068 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp 1704896540
transform 1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _086_
timestamp 1704896540
transform 1 0 46092 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp 1704896540
transform 1 0 47472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _088_
timestamp 1704896540
transform 1 0 46644 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp 1704896540
transform 1 0 49036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1704896540
transform -1 0 61364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1704896540
transform -1 0 53360 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp 1704896540
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _093_
timestamp 1704896540
transform -1 0 55016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp 1704896540
transform 1 0 54648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _095_
timestamp 1704896540
transform -1 0 56580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp 1704896540
transform 1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _097_
timestamp 1704896540
transform -1 0 58236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp 1704896540
transform 1 0 57776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _099_
timestamp 1704896540
transform -1 0 59800 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp 1704896540
transform 1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _101_
timestamp 1704896540
transform -1 0 61732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp 1704896540
transform 1 0 61180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _103_
timestamp 1704896540
transform 1 0 62928 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp 1704896540
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _105_
timestamp 1704896540
transform -1 0 65136 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _106_
timestamp 1704896540
transform -1 0 64860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _107_
timestamp 1704896540
transform 1 0 66148 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1704896540
transform -1 0 66516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _109_
timestamp 1704896540
transform -1 0 68540 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _110_
timestamp 1704896540
transform 1 0 68080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _111_
timestamp 1704896540
transform -1 0 70472 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1704896540
transform -1 0 69920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _113_
timestamp 1704896540
transform -1 0 71944 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1704896540
transform -1 0 71484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _115_
timestamp 1704896540
transform -1 0 73692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _116_
timestamp 1704896540
transform 1 0 72864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _117_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 30728 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _118_
timestamp 1704896540
transform -1 0 23736 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1704896540
transform -1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25852 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _122_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20608 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20056 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 40388 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1704896540
transform -1 0 37076 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1704896540
transform 1 0 65596 0 1 33728
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2392 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6256 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7360 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8464 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8832 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9936 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11408 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12512 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13984 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_159
timestamp 1704896540
transform 1 0 15640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1704896540
transform 1 0 18952 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_220 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21252 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21712 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1704896540
transform 1 0 24288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_337
timestamp 1704896540
transform 1 0 32016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1704896540
transform 1 0 34592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_393
timestamp 1704896540
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39468 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1704896540
transform 1 0 41952 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1704896540
transform 1 0 49680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1704896540
transform 1 0 52256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1704896540
transform 1 0 54832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1704896540
transform 1 0 57408 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_617
timestamp 1704896540
transform 1 0 57776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_642
timestamp 1704896540
transform 1 0 60076 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1704896540
transform 1 0 62560 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1704896540
transform 1 0 65136 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_707
timestamp 1704896540
transform 1 0 66056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_724
timestamp 1704896540
transform 1 0 67620 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_753
timestamp 1704896540
transform 1 0 70288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_757
timestamp 1704896540
transform 1 0 70656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_761
timestamp 1704896540
transform 1 0 71024 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1288 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2392 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3496 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4600 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6256 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7360 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8464 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9568 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10672 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11224 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11408 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12512 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13616 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14720 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15824 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16560 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21528 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_271
timestamp 1704896540
transform 1 0 25944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_297
timestamp 1704896540
transform 1 0 28336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_337
timestamp 1704896540
transform 1 0 32016 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1704896540
transform 1 0 32384 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1704896540
transform 1 0 36892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_393
timestamp 1704896540
transform 1 0 37168 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_410
timestamp 1704896540
transform 1 0 38732 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_430
timestamp 1704896540
transform 1 0 40572 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_434
timestamp 1704896540
transform 1 0 40940 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1704896540
transform 1 0 42136 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_449
timestamp 1704896540
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_454
timestamp 1704896540
transform 1 0 42780 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1704896540
transform 1 0 47288 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_505
timestamp 1704896540
transform 1 0 47472 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_509
timestamp 1704896540
transform 1 0 47840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_540
timestamp 1704896540
transform 1 0 50692 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_544
timestamp 1704896540
transform 1 0 51060 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1704896540
transform 1 0 52440 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_561
timestamp 1704896540
transform 1 0 52624 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_588
timestamp 1704896540
transform 1 0 55108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_631
timestamp 1704896540
transform 1 0 59064 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_670
timestamp 1704896540
transform 1 0 62652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_681
timestamp 1704896540
transform 1 0 63664 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_737
timestamp 1704896540
transform 1 0 68816 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_774
timestamp 1704896540
transform 1 0 72220 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_783
timestamp 1704896540
transform 1 0 73048 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_793
timestamp 1704896540
transform 1 0 73968 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3496 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8648 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 11040 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13800 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15088 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_173
timestamp 1704896540
transform 1 0 16928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 1704896540
transform 1 0 24288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_296
timestamp 1704896540
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_317
timestamp 1704896540
transform 1 0 30176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_350
timestamp 1704896540
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1704896540
transform 1 0 34316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_365
timestamp 1704896540
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_388
timestamp 1704896540
transform 1 0 36708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_400
timestamp 1704896540
transform 1 0 37812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_412
timestamp 1704896540
transform 1 0 38916 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1704896540
transform 1 0 39744 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1704896540
transform 1 0 40848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_445
timestamp 1704896540
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_449
timestamp 1704896540
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_458
timestamp 1704896540
transform 1 0 43148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_485
timestamp 1704896540
transform 1 0 45632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_489
timestamp 1704896540
transform 1 0 46000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_512
timestamp 1704896540
transform 1 0 48116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_520
timestamp 1704896540
transform 1 0 48852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_530
timestamp 1704896540
transform 1 0 49772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1704896540
transform 1 0 50048 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1704896540
transform 1 0 51152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_557
timestamp 1704896540
transform 1 0 52256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_565
timestamp 1704896540
transform 1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_576
timestamp 1704896540
transform 1 0 54004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_585
timestamp 1704896540
transform 1 0 54832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_601
timestamp 1704896540
transform 1 0 56304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_609
timestamp 1704896540
transform 1 0 57040 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_620
timestamp 1704896540
transform 1 0 58052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_632
timestamp 1704896540
transform 1 0 59156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_645
timestamp 1704896540
transform 1 0 60352 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_654
timestamp 1704896540
transform 1 0 61180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_680
timestamp 1704896540
transform 1 0 63572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_692
timestamp 1704896540
transform 1 0 64676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_701
timestamp 1704896540
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_710
timestamp 1704896540
transform 1 0 66332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_718
timestamp 1704896540
transform 1 0 67068 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_726
timestamp 1704896540
transform 1 0 67804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_738
timestamp 1704896540
transform 1 0 68908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_750
timestamp 1704896540
transform 1 0 70012 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_765
timestamp 1704896540
transform 1 0 71392 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_777
timestamp 1704896540
transform 1 0 72496 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_789
timestamp 1704896540
transform 1 0 73600 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16376 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_187
timestamp 1704896540
transform 1 0 18216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_249
timestamp 1704896540
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_261
timestamp 1704896540
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_274
timestamp 1704896540
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_295
timestamp 1704896540
transform 1 0 28152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_326
timestamp 1704896540
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 1704896540
transform 1 0 31740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_349
timestamp 1704896540
transform 1 0 33120 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_366
timestamp 1704896540
transform 1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_385
timestamp 1704896540
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1704896540
transform 1 0 37168 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1704896540
transform 1 0 38272 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1704896540
transform 1 0 39376 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1704896540
transform 1 0 40480 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1704896540
transform 1 0 41584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1704896540
transform 1 0 42136 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1704896540
transform 1 0 42320 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1704896540
transform 1 0 43424 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1704896540
transform 1 0 44528 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_485
timestamp 1704896540
transform 1 0 45632 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_491
timestamp 1704896540
transform 1 0 46184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1704896540
transform 1 0 47288 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_508
timestamp 1704896540
transform 1 0 47748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_520
timestamp 1704896540
transform 1 0 48852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_525
timestamp 1704896540
transform 1 0 49312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_537
timestamp 1704896540
transform 1 0 50416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_549
timestamp 1704896540
transform 1 0 51520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_557
timestamp 1704896540
transform 1 0 52256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_561
timestamp 1704896540
transform 1 0 52624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_567
timestamp 1704896540
transform 1 0 53176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_575
timestamp 1704896540
transform 1 0 53912 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_586
timestamp 1704896540
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_598
timestamp 1704896540
transform 1 0 56028 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_603
timestamp 1704896540
transform 1 0 56488 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1704896540
transform 1 0 57592 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_620
timestamp 1704896540
transform 1 0 58052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_632
timestamp 1704896540
transform 1 0 59156 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_638
timestamp 1704896540
transform 1 0 59708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_650
timestamp 1704896540
transform 1 0 60812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_657
timestamp 1704896540
transform 1 0 61456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_669
timestamp 1704896540
transform 1 0 62560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_673
timestamp 1704896540
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_677
timestamp 1704896540
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_689
timestamp 1704896540
transform 1 0 64400 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_694
timestamp 1704896540
transform 1 0 64860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_706
timestamp 1704896540
transform 1 0 65964 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_712
timestamp 1704896540
transform 1 0 66516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_724
timestamp 1704896540
transform 1 0 67620 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_732
timestamp 1704896540
transform 1 0 68356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_744
timestamp 1704896540
transform 1 0 69460 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_749
timestamp 1704896540
transform 1 0 69920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_761
timestamp 1704896540
transform 1 0 71024 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_766
timestamp 1704896540
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_778
timestamp 1704896540
transform 1 0 72588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1704896540
transform 1 0 73232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_797
timestamp 1704896540
transform 1 0 74336 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8648 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9936 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15088 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18952 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_217
timestamp 1704896540
transform 1 0 20976 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_229
timestamp 1704896540
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_233
timestamp 1704896540
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 1704896540
transform 1 0 23736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1704896540
transform 1 0 24104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_253
timestamp 1704896540
transform 1 0 24288 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_257
timestamp 1704896540
transform 1 0 24656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_275
timestamp 1704896540
transform 1 0 26312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_283
timestamp 1704896540
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_295
timestamp 1704896540
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1704896540
transform 1 0 29256 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1704896540
transform 1 0 29440 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_321
timestamp 1704896540
transform 1 0 30544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_327
timestamp 1704896540
transform 1 0 31096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_331
timestamp 1704896540
transform 1 0 31464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_336
timestamp 1704896540
transform 1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_342
timestamp 1704896540
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_349
timestamp 1704896540
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_361
timestamp 1704896540
transform 1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1704896540
transform 1 0 34592 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1704896540
transform 1 0 35696 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1704896540
transform 1 0 36800 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1704896540
transform 1 0 37904 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1704896540
transform 1 0 39008 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1704896540
transform 1 0 39560 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1704896540
transform 1 0 39744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1704896540
transform 1 0 40848 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1704896540
transform 1 0 41952 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1704896540
transform 1 0 43056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1704896540
transform 1 0 44160 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1704896540
transform 1 0 44712 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1704896540
transform 1 0 44896 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1704896540
transform 1 0 46000 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1704896540
transform 1 0 47104 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1704896540
transform 1 0 48208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 1704896540
transform 1 0 49312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1704896540
transform 1 0 49864 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1704896540
transform 1 0 50048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1704896540
transform 1 0 51152 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1704896540
transform 1 0 52256 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1704896540
transform 1 0 53360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1704896540
transform 1 0 54464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1704896540
transform 1 0 55016 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1704896540
transform 1 0 55200 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1704896540
transform 1 0 56304 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1704896540
transform 1 0 57408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1704896540
transform 1 0 58512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1704896540
transform 1 0 59616 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1704896540
transform 1 0 60168 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1704896540
transform 1 0 60352 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1704896540
transform 1 0 61456 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1704896540
transform 1 0 62560 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1704896540
transform 1 0 63664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1704896540
transform 1 0 64768 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1704896540
transform 1 0 65320 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1704896540
transform 1 0 65504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1704896540
transform 1 0 66608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_725
timestamp 1704896540
transform 1 0 67712 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_737
timestamp 1704896540
transform 1 0 68816 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_749
timestamp 1704896540
transform 1 0 69920 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_755
timestamp 1704896540
transform 1 0 70472 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1704896540
transform 1 0 70656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1704896540
transform 1 0 71760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1704896540
transform 1 0 72864 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_793
timestamp 1704896540
transform 1 0 73968 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6072 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10672 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11224 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13616 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16376 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_197
timestamp 1704896540
transform 1 0 19136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_204
timestamp 1704896540
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_216
timestamp 1704896540
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22816 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1704896540
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1704896540
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 26128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_287
timestamp 1704896540
transform 1 0 27416 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_294
timestamp 1704896540
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_306
timestamp 1704896540
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_320
timestamp 1704896540
transform 1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_330
timestamp 1704896540
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1704896540
transform 1 0 32016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1704896540
transform 1 0 33120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_361
timestamp 1704896540
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_365
timestamp 1704896540
transform 1 0 34592 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_370
timestamp 1704896540
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_382
timestamp 1704896540
transform 1 0 36156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1704896540
transform 1 0 36892 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1704896540
transform 1 0 37168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1704896540
transform 1 0 38272 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1704896540
transform 1 0 39376 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1704896540
transform 1 0 40480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1704896540
transform 1 0 41584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1704896540
transform 1 0 42136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1704896540
transform 1 0 42320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1704896540
transform 1 0 43424 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1704896540
transform 1 0 44528 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1704896540
transform 1 0 45632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 1704896540
transform 1 0 46736 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1704896540
transform 1 0 47288 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1704896540
transform 1 0 47472 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1704896540
transform 1 0 48576 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1704896540
transform 1 0 49680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1704896540
transform 1 0 50784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 1704896540
transform 1 0 51888 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1704896540
transform 1 0 52440 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1704896540
transform 1 0 52624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1704896540
transform 1 0 53728 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1704896540
transform 1 0 54832 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1704896540
transform 1 0 55936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1704896540
transform 1 0 57040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1704896540
transform 1 0 57592 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1704896540
transform 1 0 57776 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1704896540
transform 1 0 58880 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1704896540
transform 1 0 59984 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1704896540
transform 1 0 61088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1704896540
transform 1 0 62192 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1704896540
transform 1 0 62744 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1704896540
transform 1 0 62928 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1704896540
transform 1 0 64032 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1704896540
transform 1 0 65136 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1704896540
transform 1 0 66240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1704896540
transform 1 0 67344 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1704896540
transform 1 0 67896 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1704896540
transform 1 0 68080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1704896540
transform 1 0 69184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1704896540
transform 1 0 70288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1704896540
transform 1 0 71392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1704896540
transform 1 0 72496 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1704896540
transform 1 0 73048 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1704896540
transform 1 0 73232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_797
timestamp 1704896540
transform 1 0 74336 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8096 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8648 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9936 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13800 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15088 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23552 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 24104 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1704896540
transform 1 0 24288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1704896540
transform 1 0 25392 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1704896540
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1704896540
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1704896540
transform 1 0 28704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1704896540
transform 1 0 29256 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1704896540
transform 1 0 29440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1704896540
transform 1 0 30544 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1704896540
transform 1 0 31648 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1704896540
transform 1 0 32752 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_357
timestamp 1704896540
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1704896540
transform 1 0 34592 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1704896540
transform 1 0 35696 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1704896540
transform 1 0 36800 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1704896540
transform 1 0 37904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1704896540
transform 1 0 39008 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1704896540
transform 1 0 39560 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1704896540
transform 1 0 39744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_433
timestamp 1704896540
transform 1 0 40848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_453
timestamp 1704896540
transform 1 0 42688 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_459
timestamp 1704896540
transform 1 0 43240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_473
timestamp 1704896540
transform 1 0 44528 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1704896540
transform 1 0 44896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_489
timestamp 1704896540
transform 1 0 46000 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_495
timestamp 1704896540
transform 1 0 46552 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1704896540
transform 1 0 47104 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1704896540
transform 1 0 48208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 1704896540
transform 1 0 49312 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 1704896540
transform 1 0 49864 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1704896540
transform 1 0 50048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1704896540
transform 1 0 51152 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1704896540
transform 1 0 52256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1704896540
transform 1 0 53360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1704896540
transform 1 0 54464 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1704896540
transform 1 0 55016 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1704896540
transform 1 0 55200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1704896540
transform 1 0 56304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1704896540
transform 1 0 57408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1704896540
transform 1 0 58512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1704896540
transform 1 0 59616 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1704896540
transform 1 0 60168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_645
timestamp 1704896540
transform 1 0 60352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_651
timestamp 1704896540
transform 1 0 60904 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_656
timestamp 1704896540
transform 1 0 61364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_668
timestamp 1704896540
transform 1 0 62468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_680
timestamp 1704896540
transform 1 0 63572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_692
timestamp 1704896540
transform 1 0 64676 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1704896540
transform 1 0 65504 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1704896540
transform 1 0 66608 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1704896540
transform 1 0 67712 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1704896540
transform 1 0 68816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1704896540
transform 1 0 69920 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1704896540
transform 1 0 70472 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1704896540
transform 1 0 70656 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1704896540
transform 1 0 71760 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1704896540
transform 1 0 72864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_793
timestamp 1704896540
transform 1 0 73968 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10672 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11224 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16376 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1704896540
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1704896540
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22816 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp 1704896540
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_260
timestamp 1704896540
transform 1 0 24932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_264
timestamp 1704896540
transform 1 0 25300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_293
timestamp 1704896540
transform 1 0 27968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_299
timestamp 1704896540
transform 1 0 28520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_306
timestamp 1704896540
transform 1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_313
timestamp 1704896540
transform 1 0 29808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_319
timestamp 1704896540
transform 1 0 30360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_325
timestamp 1704896540
transform 1 0 30912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_333
timestamp 1704896540
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1704896540
transform 1 0 32016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1704896540
transform 1 0 33120 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1704896540
transform 1 0 34224 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1704896540
transform 1 0 35328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1704896540
transform 1 0 36432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1704896540
transform 1 0 36984 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1704896540
transform 1 0 37168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1704896540
transform 1 0 38272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_417
timestamp 1704896540
transform 1 0 39376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_425
timestamp 1704896540
transform 1 0 40112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_436
timestamp 1704896540
transform 1 0 41124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_449
timestamp 1704896540
transform 1 0 42320 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_455
timestamp 1704896540
transform 1 0 42872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_480
timestamp 1704896540
transform 1 0 45172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 1704896540
transform 1 0 47288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_513
timestamp 1704896540
transform 1 0 48208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_521
timestamp 1704896540
transform 1 0 48944 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_531
timestamp 1704896540
transform 1 0 49864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_543
timestamp 1704896540
transform 1 0 50968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_555
timestamp 1704896540
transform 1 0 52072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 1704896540
transform 1 0 52440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_561
timestamp 1704896540
transform 1 0 52624 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_569
timestamp 1704896540
transform 1 0 53360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_581
timestamp 1704896540
transform 1 0 54464 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_587
timestamp 1704896540
transform 1 0 55016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_599
timestamp 1704896540
transform 1 0 56120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_611
timestamp 1704896540
transform 1 0 57224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1704896540
transform 1 0 57592 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1704896540
transform 1 0 57776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1704896540
transform 1 0 58880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1704896540
transform 1 0 59984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1704896540
transform 1 0 61088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1704896540
transform 1 0 62192 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1704896540
transform 1 0 62744 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1704896540
transform 1 0 62928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1704896540
transform 1 0 64032 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1704896540
transform 1 0 65136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1704896540
transform 1 0 66240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1704896540
transform 1 0 67344 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1704896540
transform 1 0 67896 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1704896540
transform 1 0 68080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_741
timestamp 1704896540
transform 1 0 69184 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_749
timestamp 1704896540
transform 1 0 69920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_755
timestamp 1704896540
transform 1 0 70472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_763
timestamp 1704896540
transform 1 0 71208 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_771
timestamp 1704896540
transform 1 0 71944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1704896540
transform 1 0 73048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_790
timestamp 1704896540
transform 1 0 73692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_798
timestamp 1704896540
transform 1 0 74428 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1704896540
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1704896540
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1704896540
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_113
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1704896540
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1704896540
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_169
timestamp 1704896540
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_181
timestamp 1704896540
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1704896540
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 20240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_221
timestamp 1704896540
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_225
timestamp 1704896540
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_237
timestamp 1704896540
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_241
timestamp 1704896540
transform 1 0 23184 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_263
timestamp 1704896540
transform 1 0 25208 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_274
timestamp 1704896540
transform 1 0 26220 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_281
timestamp 1704896540
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_293
timestamp 1704896540
transform 1 0 27968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 1704896540
transform 1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1704896540
transform 1 0 29440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1704896540
transform 1 0 30544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_333
timestamp 1704896540
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_337
timestamp 1704896540
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_349
timestamp 1704896540
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1704896540
transform 1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_365
timestamp 1704896540
transform 1 0 34592 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_371
timestamp 1704896540
transform 1 0 35144 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_393
timestamp 1704896540
transform 1 0 37168 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_405
timestamp 1704896540
transform 1 0 38272 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_417
timestamp 1704896540
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_421
timestamp 1704896540
transform 1 0 39744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_427
timestamp 1704896540
transform 1 0 40296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1704896540
transform 1 0 44528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_501
timestamp 1704896540
transform 1 0 47104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_529
timestamp 1704896540
transform 1 0 49680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_533
timestamp 1704896540
transform 1 0 50048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_545
timestamp 1704896540
transform 1 0 51152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_554
timestamp 1704896540
transform 1 0 51980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_585
timestamp 1704896540
transform 1 0 54832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_597
timestamp 1704896540
transform 1 0 55936 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_604
timestamp 1704896540
transform 1 0 56580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_622
timestamp 1704896540
transform 1 0 58236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_639
timestamp 1704896540
transform 1 0 59800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1704896540
transform 1 0 60168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_645
timestamp 1704896540
transform 1 0 60352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_653
timestamp 1704896540
transform 1 0 61088 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_660
timestamp 1704896540
transform 1 0 61732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_678
timestamp 1704896540
transform 1 0 63388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_690
timestamp 1704896540
transform 1 0 64492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_697
timestamp 1704896540
transform 1 0 65136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_701
timestamp 1704896540
transform 1 0 65504 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_707
timestamp 1704896540
transform 1 0 66056 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1704896540
transform 1 0 66608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_725
timestamp 1704896540
transform 1 0 67712 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_734
timestamp 1704896540
transform 1 0 68540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_746
timestamp 1704896540
transform 1 0 69644 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_754
timestamp 1704896540
transform 1 0 70380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1704896540
transform 1 0 70656 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1704896540
transform 1 0 71760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_781
timestamp 1704896540
transform 1 0 72864 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_785
timestamp 1704896540
transform 1 0 73232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_797
timestamp 1704896540
transform 1 0 74336 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_702
timestamp 1704896540
transform 1 0 65596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_714
timestamp 1704896540
transform 1 0 66700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_726
timestamp 1704896540
transform 1 0 67804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_738
timestamp 1704896540
transform 1 0 68908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_750
timestamp 1704896540
transform 1 0 70012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_754
timestamp 1704896540
transform 1 0 70380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_756
timestamp 1704896540
transform 1 0 70564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_768
timestamp 1704896540
transform 1 0 71668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_780
timestamp 1704896540
transform 1 0 72772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_792
timestamp 1704896540
transform 1 0 73876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_800
timestamp 1704896540
transform 1 0 74612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_702
timestamp 1704896540
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_714
timestamp 1704896540
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_726
timestamp 1704896540
transform 1 0 67804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_728
timestamp 1704896540
transform 1 0 67988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_740
timestamp 1704896540
transform 1 0 69092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_752
timestamp 1704896540
transform 1 0 70196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_764
timestamp 1704896540
transform 1 0 71300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_776
timestamp 1704896540
transform 1 0 72404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_782
timestamp 1704896540
transform 1 0 72956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_784
timestamp 1704896540
transform 1 0 73140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_796
timestamp 1704896540
transform 1 0 74244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_800
timestamp 1704896540
transform 1 0 74612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_702
timestamp 1704896540
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_714
timestamp 1704896540
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_726
timestamp 1704896540
transform 1 0 67804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_738
timestamp 1704896540
transform 1 0 68908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_750
timestamp 1704896540
transform 1 0 70012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_754
timestamp 1704896540
transform 1 0 70380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_756
timestamp 1704896540
transform 1 0 70564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_768
timestamp 1704896540
transform 1 0 71668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_780
timestamp 1704896540
transform 1 0 72772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_792
timestamp 1704896540
transform 1 0 73876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_800
timestamp 1704896540
transform 1 0 74612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_702
timestamp 1704896540
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_714
timestamp 1704896540
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_726
timestamp 1704896540
transform 1 0 67804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_728
timestamp 1704896540
transform 1 0 67988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_740
timestamp 1704896540
transform 1 0 69092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_752
timestamp 1704896540
transform 1 0 70196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_764
timestamp 1704896540
transform 1 0 71300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_776
timestamp 1704896540
transform 1 0 72404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_782
timestamp 1704896540
transform 1 0 72956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_784
timestamp 1704896540
transform 1 0 73140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_796
timestamp 1704896540
transform 1 0 74244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_800
timestamp 1704896540
transform 1 0 74612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_702
timestamp 1704896540
transform 1 0 65596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_714
timestamp 1704896540
transform 1 0 66700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_726
timestamp 1704896540
transform 1 0 67804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_738
timestamp 1704896540
transform 1 0 68908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_750
timestamp 1704896540
transform 1 0 70012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_754
timestamp 1704896540
transform 1 0 70380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_756
timestamp 1704896540
transform 1 0 70564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_768
timestamp 1704896540
transform 1 0 71668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_780
timestamp 1704896540
transform 1 0 72772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_792
timestamp 1704896540
transform 1 0 73876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_800
timestamp 1704896540
transform 1 0 74612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_702
timestamp 1704896540
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_714
timestamp 1704896540
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_726
timestamp 1704896540
transform 1 0 67804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_728
timestamp 1704896540
transform 1 0 67988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_740
timestamp 1704896540
transform 1 0 69092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_752
timestamp 1704896540
transform 1 0 70196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_764
timestamp 1704896540
transform 1 0 71300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_776
timestamp 1704896540
transform 1 0 72404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_782
timestamp 1704896540
transform 1 0 72956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_784
timestamp 1704896540
transform 1 0 73140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_796
timestamp 1704896540
transform 1 0 74244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_800
timestamp 1704896540
transform 1 0 74612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_702
timestamp 1704896540
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_714
timestamp 1704896540
transform 1 0 66700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_726
timestamp 1704896540
transform 1 0 67804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_738
timestamp 1704896540
transform 1 0 68908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_750
timestamp 1704896540
transform 1 0 70012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_754
timestamp 1704896540
transform 1 0 70380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_756
timestamp 1704896540
transform 1 0 70564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_768
timestamp 1704896540
transform 1 0 71668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_780
timestamp 1704896540
transform 1 0 72772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_792
timestamp 1704896540
transform 1 0 73876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_800
timestamp 1704896540
transform 1 0 74612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_702
timestamp 1704896540
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_714
timestamp 1704896540
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_726
timestamp 1704896540
transform 1 0 67804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_728
timestamp 1704896540
transform 1 0 67988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_740
timestamp 1704896540
transform 1 0 69092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_752
timestamp 1704896540
transform 1 0 70196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_764
timestamp 1704896540
transform 1 0 71300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_776
timestamp 1704896540
transform 1 0 72404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_782
timestamp 1704896540
transform 1 0 72956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_784
timestamp 1704896540
transform 1 0 73140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_796
timestamp 1704896540
transform 1 0 74244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_800
timestamp 1704896540
transform 1 0 74612 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_702
timestamp 1704896540
transform 1 0 65596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_714
timestamp 1704896540
transform 1 0 66700 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_726
timestamp 1704896540
transform 1 0 67804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_738
timestamp 1704896540
transform 1 0 68908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_750
timestamp 1704896540
transform 1 0 70012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_754
timestamp 1704896540
transform 1 0 70380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_756
timestamp 1704896540
transform 1 0 70564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_768
timestamp 1704896540
transform 1 0 71668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_780
timestamp 1704896540
transform 1 0 72772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_792
timestamp 1704896540
transform 1 0 73876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_800
timestamp 1704896540
transform 1 0 74612 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_702
timestamp 1704896540
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_714
timestamp 1704896540
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_726
timestamp 1704896540
transform 1 0 67804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_728
timestamp 1704896540
transform 1 0 67988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_740
timestamp 1704896540
transform 1 0 69092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_752
timestamp 1704896540
transform 1 0 70196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_764
timestamp 1704896540
transform 1 0 71300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_776
timestamp 1704896540
transform 1 0 72404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_782
timestamp 1704896540
transform 1 0 72956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_784
timestamp 1704896540
transform 1 0 73140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_796
timestamp 1704896540
transform 1 0 74244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_800
timestamp 1704896540
transform 1 0 74612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_702
timestamp 1704896540
transform 1 0 65596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_714
timestamp 1704896540
transform 1 0 66700 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_726
timestamp 1704896540
transform 1 0 67804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_738
timestamp 1704896540
transform 1 0 68908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_750
timestamp 1704896540
transform 1 0 70012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_754
timestamp 1704896540
transform 1 0 70380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_756
timestamp 1704896540
transform 1 0 70564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_768
timestamp 1704896540
transform 1 0 71668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_780
timestamp 1704896540
transform 1 0 72772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_792
timestamp 1704896540
transform 1 0 73876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_800
timestamp 1704896540
transform 1 0 74612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_702
timestamp 1704896540
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_714
timestamp 1704896540
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_726
timestamp 1704896540
transform 1 0 67804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_728
timestamp 1704896540
transform 1 0 67988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_740
timestamp 1704896540
transform 1 0 69092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_752
timestamp 1704896540
transform 1 0 70196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_764
timestamp 1704896540
transform 1 0 71300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_776
timestamp 1704896540
transform 1 0 72404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_782
timestamp 1704896540
transform 1 0 72956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_784
timestamp 1704896540
transform 1 0 73140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_796
timestamp 1704896540
transform 1 0 74244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_800
timestamp 1704896540
transform 1 0 74612 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_702
timestamp 1704896540
transform 1 0 65596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_714
timestamp 1704896540
transform 1 0 66700 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_726
timestamp 1704896540
transform 1 0 67804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_738
timestamp 1704896540
transform 1 0 68908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_750
timestamp 1704896540
transform 1 0 70012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_754
timestamp 1704896540
transform 1 0 70380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_756
timestamp 1704896540
transform 1 0 70564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_768
timestamp 1704896540
transform 1 0 71668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_780
timestamp 1704896540
transform 1 0 72772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_792
timestamp 1704896540
transform 1 0 73876 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_800
timestamp 1704896540
transform 1 0 74612 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_702
timestamp 1704896540
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_714
timestamp 1704896540
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_726
timestamp 1704896540
transform 1 0 67804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_728
timestamp 1704896540
transform 1 0 67988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_740
timestamp 1704896540
transform 1 0 69092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_752
timestamp 1704896540
transform 1 0 70196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_764
timestamp 1704896540
transform 1 0 71300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_776
timestamp 1704896540
transform 1 0 72404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_782
timestamp 1704896540
transform 1 0 72956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_784
timestamp 1704896540
transform 1 0 73140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_796
timestamp 1704896540
transform 1 0 74244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_800
timestamp 1704896540
transform 1 0 74612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_702
timestamp 1704896540
transform 1 0 65596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_714
timestamp 1704896540
transform 1 0 66700 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_726
timestamp 1704896540
transform 1 0 67804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_738
timestamp 1704896540
transform 1 0 68908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_750
timestamp 1704896540
transform 1 0 70012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_754
timestamp 1704896540
transform 1 0 70380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_756
timestamp 1704896540
transform 1 0 70564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_768
timestamp 1704896540
transform 1 0 71668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_780
timestamp 1704896540
transform 1 0 72772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_792
timestamp 1704896540
transform 1 0 73876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_800
timestamp 1704896540
transform 1 0 74612 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_702
timestamp 1704896540
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_714
timestamp 1704896540
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_726
timestamp 1704896540
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_728
timestamp 1704896540
transform 1 0 67988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_740
timestamp 1704896540
transform 1 0 69092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_752
timestamp 1704896540
transform 1 0 70196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_764
timestamp 1704896540
transform 1 0 71300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_776
timestamp 1704896540
transform 1 0 72404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_782
timestamp 1704896540
transform 1 0 72956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_784
timestamp 1704896540
transform 1 0 73140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_796
timestamp 1704896540
transform 1 0 74244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_800
timestamp 1704896540
transform 1 0 74612 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_702
timestamp 1704896540
transform 1 0 65596 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_714
timestamp 1704896540
transform 1 0 66700 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_726
timestamp 1704896540
transform 1 0 67804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_738
timestamp 1704896540
transform 1 0 68908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_750
timestamp 1704896540
transform 1 0 70012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_754
timestamp 1704896540
transform 1 0 70380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_756
timestamp 1704896540
transform 1 0 70564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_768
timestamp 1704896540
transform 1 0 71668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_780
timestamp 1704896540
transform 1 0 72772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_792
timestamp 1704896540
transform 1 0 73876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_800
timestamp 1704896540
transform 1 0 74612 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_702
timestamp 1704896540
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_714
timestamp 1704896540
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_726
timestamp 1704896540
transform 1 0 67804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_728
timestamp 1704896540
transform 1 0 67988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_740
timestamp 1704896540
transform 1 0 69092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_752
timestamp 1704896540
transform 1 0 70196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_764
timestamp 1704896540
transform 1 0 71300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_776
timestamp 1704896540
transform 1 0 72404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_782
timestamp 1704896540
transform 1 0 72956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_784
timestamp 1704896540
transform 1 0 73140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_796
timestamp 1704896540
transform 1 0 74244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_800
timestamp 1704896540
transform 1 0 74612 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_702
timestamp 1704896540
transform 1 0 65596 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_714
timestamp 1704896540
transform 1 0 66700 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_726
timestamp 1704896540
transform 1 0 67804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_738
timestamp 1704896540
transform 1 0 68908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_750
timestamp 1704896540
transform 1 0 70012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_754
timestamp 1704896540
transform 1 0 70380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_756
timestamp 1704896540
transform 1 0 70564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_768
timestamp 1704896540
transform 1 0 71668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_780
timestamp 1704896540
transform 1 0 72772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_792
timestamp 1704896540
transform 1 0 73876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_800
timestamp 1704896540
transform 1 0 74612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_702
timestamp 1704896540
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_714
timestamp 1704896540
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_726
timestamp 1704896540
transform 1 0 67804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_728
timestamp 1704896540
transform 1 0 67988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_740
timestamp 1704896540
transform 1 0 69092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_752
timestamp 1704896540
transform 1 0 70196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_764
timestamp 1704896540
transform 1 0 71300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_776
timestamp 1704896540
transform 1 0 72404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_782
timestamp 1704896540
transform 1 0 72956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_784
timestamp 1704896540
transform 1 0 73140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_796
timestamp 1704896540
transform 1 0 74244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_800
timestamp 1704896540
transform 1 0 74612 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_702
timestamp 1704896540
transform 1 0 65596 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_714
timestamp 1704896540
transform 1 0 66700 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_726
timestamp 1704896540
transform 1 0 67804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_738
timestamp 1704896540
transform 1 0 68908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_750
timestamp 1704896540
transform 1 0 70012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_754
timestamp 1704896540
transform 1 0 70380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_756
timestamp 1704896540
transform 1 0 70564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_768
timestamp 1704896540
transform 1 0 71668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_780
timestamp 1704896540
transform 1 0 72772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_792
timestamp 1704896540
transform 1 0 73876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_800
timestamp 1704896540
transform 1 0 74612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_702
timestamp 1704896540
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_714
timestamp 1704896540
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_726
timestamp 1704896540
transform 1 0 67804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_728
timestamp 1704896540
transform 1 0 67988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_740
timestamp 1704896540
transform 1 0 69092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_752
timestamp 1704896540
transform 1 0 70196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_764
timestamp 1704896540
transform 1 0 71300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_776
timestamp 1704896540
transform 1 0 72404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_782
timestamp 1704896540
transform 1 0 72956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_784
timestamp 1704896540
transform 1 0 73140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_796
timestamp 1704896540
transform 1 0 74244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_800
timestamp 1704896540
transform 1 0 74612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_702
timestamp 1704896540
transform 1 0 65596 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_714
timestamp 1704896540
transform 1 0 66700 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_726
timestamp 1704896540
transform 1 0 67804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_738
timestamp 1704896540
transform 1 0 68908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_750
timestamp 1704896540
transform 1 0 70012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_754
timestamp 1704896540
transform 1 0 70380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_756
timestamp 1704896540
transform 1 0 70564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_768
timestamp 1704896540
transform 1 0 71668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_780
timestamp 1704896540
transform 1 0 72772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_792
timestamp 1704896540
transform 1 0 73876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_800
timestamp 1704896540
transform 1 0 74612 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_702
timestamp 1704896540
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_714
timestamp 1704896540
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_726
timestamp 1704896540
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_728
timestamp 1704896540
transform 1 0 67988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_740
timestamp 1704896540
transform 1 0 69092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_752
timestamp 1704896540
transform 1 0 70196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_764
timestamp 1704896540
transform 1 0 71300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_776
timestamp 1704896540
transform 1 0 72404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_782
timestamp 1704896540
transform 1 0 72956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_784
timestamp 1704896540
transform 1 0 73140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_796
timestamp 1704896540
transform 1 0 74244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_800
timestamp 1704896540
transform 1 0 74612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_702
timestamp 1704896540
transform 1 0 65596 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_714
timestamp 1704896540
transform 1 0 66700 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_726
timestamp 1704896540
transform 1 0 67804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_738
timestamp 1704896540
transform 1 0 68908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_750
timestamp 1704896540
transform 1 0 70012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_754
timestamp 1704896540
transform 1 0 70380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_756
timestamp 1704896540
transform 1 0 70564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_768
timestamp 1704896540
transform 1 0 71668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_780
timestamp 1704896540
transform 1 0 72772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_792
timestamp 1704896540
transform 1 0 73876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_800
timestamp 1704896540
transform 1 0 74612 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_702
timestamp 1704896540
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_714
timestamp 1704896540
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_726
timestamp 1704896540
transform 1 0 67804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_728
timestamp 1704896540
transform 1 0 67988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_740
timestamp 1704896540
transform 1 0 69092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_752
timestamp 1704896540
transform 1 0 70196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_764
timestamp 1704896540
transform 1 0 71300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_776
timestamp 1704896540
transform 1 0 72404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_782
timestamp 1704896540
transform 1 0 72956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_784
timestamp 1704896540
transform 1 0 73140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_796
timestamp 1704896540
transform 1 0 74244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_800
timestamp 1704896540
transform 1 0 74612 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_702
timestamp 1704896540
transform 1 0 65596 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_714
timestamp 1704896540
transform 1 0 66700 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_726
timestamp 1704896540
transform 1 0 67804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_738
timestamp 1704896540
transform 1 0 68908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_750
timestamp 1704896540
transform 1 0 70012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_754
timestamp 1704896540
transform 1 0 70380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_756
timestamp 1704896540
transform 1 0 70564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_768
timestamp 1704896540
transform 1 0 71668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_780
timestamp 1704896540
transform 1 0 72772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_792
timestamp 1704896540
transform 1 0 73876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_800
timestamp 1704896540
transform 1 0 74612 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_702
timestamp 1704896540
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_714
timestamp 1704896540
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_726
timestamp 1704896540
transform 1 0 67804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_728
timestamp 1704896540
transform 1 0 67988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_740
timestamp 1704896540
transform 1 0 69092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_752
timestamp 1704896540
transform 1 0 70196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_764
timestamp 1704896540
transform 1 0 71300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_776
timestamp 1704896540
transform 1 0 72404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_782
timestamp 1704896540
transform 1 0 72956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_784
timestamp 1704896540
transform 1 0 73140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_796
timestamp 1704896540
transform 1 0 74244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_800
timestamp 1704896540
transform 1 0 74612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_702
timestamp 1704896540
transform 1 0 65596 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_714
timestamp 1704896540
transform 1 0 66700 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_726
timestamp 1704896540
transform 1 0 67804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_738
timestamp 1704896540
transform 1 0 68908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_750
timestamp 1704896540
transform 1 0 70012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_754
timestamp 1704896540
transform 1 0 70380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_756
timestamp 1704896540
transform 1 0 70564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_768
timestamp 1704896540
transform 1 0 71668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_780
timestamp 1704896540
transform 1 0 72772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_792
timestamp 1704896540
transform 1 0 73876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_800
timestamp 1704896540
transform 1 0 74612 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_702
timestamp 1704896540
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_714
timestamp 1704896540
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_726
timestamp 1704896540
transform 1 0 67804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_728
timestamp 1704896540
transform 1 0 67988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_740
timestamp 1704896540
transform 1 0 69092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_752
timestamp 1704896540
transform 1 0 70196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_764
timestamp 1704896540
transform 1 0 71300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_776
timestamp 1704896540
transform 1 0 72404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_782
timestamp 1704896540
transform 1 0 72956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_784
timestamp 1704896540
transform 1 0 73140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_796
timestamp 1704896540
transform 1 0 74244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_800
timestamp 1704896540
transform 1 0 74612 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_702
timestamp 1704896540
transform 1 0 65596 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_714
timestamp 1704896540
transform 1 0 66700 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_726
timestamp 1704896540
transform 1 0 67804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_738
timestamp 1704896540
transform 1 0 68908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_750
timestamp 1704896540
transform 1 0 70012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_754
timestamp 1704896540
transform 1 0 70380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_756
timestamp 1704896540
transform 1 0 70564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_768
timestamp 1704896540
transform 1 0 71668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_780
timestamp 1704896540
transform 1 0 72772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_792
timestamp 1704896540
transform 1 0 73876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_800
timestamp 1704896540
transform 1 0 74612 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_710
timestamp 1704896540
transform 1 0 66332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_722
timestamp 1704896540
transform 1 0 67436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_726
timestamp 1704896540
transform 1 0 67804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_728
timestamp 1704896540
transform 1 0 67988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_740
timestamp 1704896540
transform 1 0 69092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_752
timestamp 1704896540
transform 1 0 70196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_764
timestamp 1704896540
transform 1 0 71300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_776
timestamp 1704896540
transform 1 0 72404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_782
timestamp 1704896540
transform 1 0 72956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_784
timestamp 1704896540
transform 1 0 73140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_796
timestamp 1704896540
transform 1 0 74244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_800
timestamp 1704896540
transform 1 0 74612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_710
timestamp 1704896540
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_722
timestamp 1704896540
transform 1 0 67436 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_734
timestamp 1704896540
transform 1 0 68540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_746
timestamp 1704896540
transform 1 0 69644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_754
timestamp 1704896540
transform 1 0 70380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_756
timestamp 1704896540
transform 1 0 70564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_768
timestamp 1704896540
transform 1 0 71668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_780
timestamp 1704896540
transform 1 0 72772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_792
timestamp 1704896540
transform 1 0 73876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_800
timestamp 1704896540
transform 1 0 74612 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_710
timestamp 1704896540
transform 1 0 66332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_722
timestamp 1704896540
transform 1 0 67436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_726
timestamp 1704896540
transform 1 0 67804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_728
timestamp 1704896540
transform 1 0 67988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_740
timestamp 1704896540
transform 1 0 69092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_752
timestamp 1704896540
transform 1 0 70196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_764
timestamp 1704896540
transform 1 0 71300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_776
timestamp 1704896540
transform 1 0 72404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_782
timestamp 1704896540
transform 1 0 72956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_784
timestamp 1704896540
transform 1 0 73140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_796
timestamp 1704896540
transform 1 0 74244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_800
timestamp 1704896540
transform 1 0 74612 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_702
timestamp 1704896540
transform 1 0 65596 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_714
timestamp 1704896540
transform 1 0 66700 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_726
timestamp 1704896540
transform 1 0 67804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_738
timestamp 1704896540
transform 1 0 68908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_750
timestamp 1704896540
transform 1 0 70012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_754
timestamp 1704896540
transform 1 0 70380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_756
timestamp 1704896540
transform 1 0 70564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_768
timestamp 1704896540
transform 1 0 71668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_780
timestamp 1704896540
transform 1 0 72772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_792
timestamp 1704896540
transform 1 0 73876 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_800
timestamp 1704896540
transform 1 0 74612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_702
timestamp 1704896540
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_714
timestamp 1704896540
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_726
timestamp 1704896540
transform 1 0 67804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_728
timestamp 1704896540
transform 1 0 67988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_740
timestamp 1704896540
transform 1 0 69092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_752
timestamp 1704896540
transform 1 0 70196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_764
timestamp 1704896540
transform 1 0 71300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_776
timestamp 1704896540
transform 1 0 72404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_782
timestamp 1704896540
transform 1 0 72956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_784
timestamp 1704896540
transform 1 0 73140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_796
timestamp 1704896540
transform 1 0 74244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_800
timestamp 1704896540
transform 1 0 74612 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_702
timestamp 1704896540
transform 1 0 65596 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_714
timestamp 1704896540
transform 1 0 66700 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_726
timestamp 1704896540
transform 1 0 67804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_738
timestamp 1704896540
transform 1 0 68908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_750
timestamp 1704896540
transform 1 0 70012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_754
timestamp 1704896540
transform 1 0 70380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_756
timestamp 1704896540
transform 1 0 70564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_768
timestamp 1704896540
transform 1 0 71668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_780
timestamp 1704896540
transform 1 0 72772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_792
timestamp 1704896540
transform 1 0 73876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_800
timestamp 1704896540
transform 1 0 74612 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_710
timestamp 1704896540
transform 1 0 66332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_722
timestamp 1704896540
transform 1 0 67436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_726
timestamp 1704896540
transform 1 0 67804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_728
timestamp 1704896540
transform 1 0 67988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_740
timestamp 1704896540
transform 1 0 69092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_752
timestamp 1704896540
transform 1 0 70196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_764
timestamp 1704896540
transform 1 0 71300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_776
timestamp 1704896540
transform 1 0 72404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_782
timestamp 1704896540
transform 1 0 72956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_784
timestamp 1704896540
transform 1 0 73140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_796
timestamp 1704896540
transform 1 0 74244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_800
timestamp 1704896540
transform 1 0 74612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_718
timestamp 1704896540
transform 1 0 67068 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_730
timestamp 1704896540
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_742
timestamp 1704896540
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_754
timestamp 1704896540
transform 1 0 70380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_756
timestamp 1704896540
transform 1 0 70564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_768
timestamp 1704896540
transform 1 0 71668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_780
timestamp 1704896540
transform 1 0 72772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_792
timestamp 1704896540
transform 1 0 73876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_800
timestamp 1704896540
transform 1 0 74612 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_710
timestamp 1704896540
transform 1 0 66332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_722
timestamp 1704896540
transform 1 0 67436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_726
timestamp 1704896540
transform 1 0 67804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_728
timestamp 1704896540
transform 1 0 67988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_740
timestamp 1704896540
transform 1 0 69092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_752
timestamp 1704896540
transform 1 0 70196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_764
timestamp 1704896540
transform 1 0 71300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_776
timestamp 1704896540
transform 1 0 72404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_782
timestamp 1704896540
transform 1 0 72956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_784
timestamp 1704896540
transform 1 0 73140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_796
timestamp 1704896540
transform 1 0 74244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_800
timestamp 1704896540
transform 1 0 74612 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_702
timestamp 1704896540
transform 1 0 65596 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_714
timestamp 1704896540
transform 1 0 66700 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_726
timestamp 1704896540
transform 1 0 67804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_738
timestamp 1704896540
transform 1 0 68908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_750
timestamp 1704896540
transform 1 0 70012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_754
timestamp 1704896540
transform 1 0 70380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_756
timestamp 1704896540
transform 1 0 70564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_768
timestamp 1704896540
transform 1 0 71668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_780
timestamp 1704896540
transform 1 0 72772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_792
timestamp 1704896540
transform 1 0 73876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_800
timestamp 1704896540
transform 1 0 74612 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_710
timestamp 1704896540
transform 1 0 66332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_722
timestamp 1704896540
transform 1 0 67436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_726
timestamp 1704896540
transform 1 0 67804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_728
timestamp 1704896540
transform 1 0 67988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_740
timestamp 1704896540
transform 1 0 69092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_752
timestamp 1704896540
transform 1 0 70196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_764
timestamp 1704896540
transform 1 0 71300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_776
timestamp 1704896540
transform 1 0 72404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_782
timestamp 1704896540
transform 1 0 72956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_784
timestamp 1704896540
transform 1 0 73140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_796
timestamp 1704896540
transform 1 0 74244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_800
timestamp 1704896540
transform 1 0 74612 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_702
timestamp 1704896540
transform 1 0 65596 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_714
timestamp 1704896540
transform 1 0 66700 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_726
timestamp 1704896540
transform 1 0 67804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_738
timestamp 1704896540
transform 1 0 68908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_750
timestamp 1704896540
transform 1 0 70012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_754
timestamp 1704896540
transform 1 0 70380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_756
timestamp 1704896540
transform 1 0 70564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_768
timestamp 1704896540
transform 1 0 71668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_780
timestamp 1704896540
transform 1 0 72772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_792
timestamp 1704896540
transform 1 0 73876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_800
timestamp 1704896540
transform 1 0 74612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_710
timestamp 1704896540
transform 1 0 66332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_722
timestamp 1704896540
transform 1 0 67436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_726
timestamp 1704896540
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_728
timestamp 1704896540
transform 1 0 67988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_740
timestamp 1704896540
transform 1 0 69092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_752
timestamp 1704896540
transform 1 0 70196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_764
timestamp 1704896540
transform 1 0 71300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_776
timestamp 1704896540
transform 1 0 72404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_782
timestamp 1704896540
transform 1 0 72956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_784
timestamp 1704896540
transform 1 0 73140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_796
timestamp 1704896540
transform 1 0 74244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_800
timestamp 1704896540
transform 1 0 74612 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_702
timestamp 1704896540
transform 1 0 65596 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_714
timestamp 1704896540
transform 1 0 66700 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_726
timestamp 1704896540
transform 1 0 67804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_738
timestamp 1704896540
transform 1 0 68908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_750
timestamp 1704896540
transform 1 0 70012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_754
timestamp 1704896540
transform 1 0 70380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_756
timestamp 1704896540
transform 1 0 70564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_768
timestamp 1704896540
transform 1 0 71668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_780
timestamp 1704896540
transform 1 0 72772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_792
timestamp 1704896540
transform 1 0 73876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_800
timestamp 1704896540
transform 1 0 74612 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_710
timestamp 1704896540
transform 1 0 66332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_722
timestamp 1704896540
transform 1 0 67436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_726
timestamp 1704896540
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_728
timestamp 1704896540
transform 1 0 67988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_740
timestamp 1704896540
transform 1 0 69092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_752
timestamp 1704896540
transform 1 0 70196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_764
timestamp 1704896540
transform 1 0 71300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_776
timestamp 1704896540
transform 1 0 72404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_782
timestamp 1704896540
transform 1 0 72956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_784
timestamp 1704896540
transform 1 0 73140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_796
timestamp 1704896540
transform 1 0 74244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_800
timestamp 1704896540
transform 1 0 74612 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_702
timestamp 1704896540
transform 1 0 65596 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_714
timestamp 1704896540
transform 1 0 66700 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_726
timestamp 1704896540
transform 1 0 67804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_738
timestamp 1704896540
transform 1 0 68908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_750
timestamp 1704896540
transform 1 0 70012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_754
timestamp 1704896540
transform 1 0 70380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_756
timestamp 1704896540
transform 1 0 70564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_768
timestamp 1704896540
transform 1 0 71668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_780
timestamp 1704896540
transform 1 0 72772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_792
timestamp 1704896540
transform 1 0 73876 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_800
timestamp 1704896540
transform 1 0 74612 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_710
timestamp 1704896540
transform 1 0 66332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_722
timestamp 1704896540
transform 1 0 67436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_726
timestamp 1704896540
transform 1 0 67804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_728
timestamp 1704896540
transform 1 0 67988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_740
timestamp 1704896540
transform 1 0 69092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_752
timestamp 1704896540
transform 1 0 70196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_764
timestamp 1704896540
transform 1 0 71300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_776
timestamp 1704896540
transform 1 0 72404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_782
timestamp 1704896540
transform 1 0 72956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_784
timestamp 1704896540
transform 1 0 73140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_796
timestamp 1704896540
transform 1 0 74244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_800
timestamp 1704896540
transform 1 0 74612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_702
timestamp 1704896540
transform 1 0 65596 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_714
timestamp 1704896540
transform 1 0 66700 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_726
timestamp 1704896540
transform 1 0 67804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_738
timestamp 1704896540
transform 1 0 68908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_750
timestamp 1704896540
transform 1 0 70012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_754
timestamp 1704896540
transform 1 0 70380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_756
timestamp 1704896540
transform 1 0 70564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_768
timestamp 1704896540
transform 1 0 71668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_780
timestamp 1704896540
transform 1 0 72772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_792
timestamp 1704896540
transform 1 0 73876 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_800
timestamp 1704896540
transform 1 0 74612 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_710
timestamp 1704896540
transform 1 0 66332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_722
timestamp 1704896540
transform 1 0 67436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_726
timestamp 1704896540
transform 1 0 67804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_728
timestamp 1704896540
transform 1 0 67988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_740
timestamp 1704896540
transform 1 0 69092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_752
timestamp 1704896540
transform 1 0 70196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_764
timestamp 1704896540
transform 1 0 71300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_776
timestamp 1704896540
transform 1 0 72404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_782
timestamp 1704896540
transform 1 0 72956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_784
timestamp 1704896540
transform 1 0 73140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_796
timestamp 1704896540
transform 1 0 74244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_800
timestamp 1704896540
transform 1 0 74612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_710
timestamp 1704896540
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_722
timestamp 1704896540
transform 1 0 67436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_734
timestamp 1704896540
transform 1 0 68540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_746
timestamp 1704896540
transform 1 0 69644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_754
timestamp 1704896540
transform 1 0 70380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_756
timestamp 1704896540
transform 1 0 70564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_768
timestamp 1704896540
transform 1 0 71668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_780
timestamp 1704896540
transform 1 0 72772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_792
timestamp 1704896540
transform 1 0 73876 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_800
timestamp 1704896540
transform 1 0 74612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_722
timestamp 1704896540
transform 1 0 67436 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_726
timestamp 1704896540
transform 1 0 67804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_728
timestamp 1704896540
transform 1 0 67988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_740
timestamp 1704896540
transform 1 0 69092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_752
timestamp 1704896540
transform 1 0 70196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_764
timestamp 1704896540
transform 1 0 71300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_776
timestamp 1704896540
transform 1 0 72404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_782
timestamp 1704896540
transform 1 0 72956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_784
timestamp 1704896540
transform 1 0 73140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_796
timestamp 1704896540
transform 1 0 74244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_800
timestamp 1704896540
transform 1 0 74612 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_702
timestamp 1704896540
transform 1 0 65596 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_714
timestamp 1704896540
transform 1 0 66700 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_726
timestamp 1704896540
transform 1 0 67804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_738
timestamp 1704896540
transform 1 0 68908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_750
timestamp 1704896540
transform 1 0 70012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_754
timestamp 1704896540
transform 1 0 70380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_756
timestamp 1704896540
transform 1 0 70564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_768
timestamp 1704896540
transform 1 0 71668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_780
timestamp 1704896540
transform 1 0 72772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_792
timestamp 1704896540
transform 1 0 73876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_800
timestamp 1704896540
transform 1 0 74612 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_710
timestamp 1704896540
transform 1 0 66332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_722
timestamp 1704896540
transform 1 0 67436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_726
timestamp 1704896540
transform 1 0 67804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_728
timestamp 1704896540
transform 1 0 67988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_740
timestamp 1704896540
transform 1 0 69092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_752
timestamp 1704896540
transform 1 0 70196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_764
timestamp 1704896540
transform 1 0 71300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_776
timestamp 1704896540
transform 1 0 72404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_782
timestamp 1704896540
transform 1 0 72956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_784
timestamp 1704896540
transform 1 0 73140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_796
timestamp 1704896540
transform 1 0 74244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_800
timestamp 1704896540
transform 1 0 74612 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_718
timestamp 1704896540
transform 1 0 67068 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_730
timestamp 1704896540
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_742
timestamp 1704896540
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_754
timestamp 1704896540
transform 1 0 70380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_756
timestamp 1704896540
transform 1 0 70564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_768
timestamp 1704896540
transform 1 0 71668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_780
timestamp 1704896540
transform 1 0 72772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_792
timestamp 1704896540
transform 1 0 73876 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_800
timestamp 1704896540
transform 1 0 74612 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_710
timestamp 1704896540
transform 1 0 66332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_722
timestamp 1704896540
transform 1 0 67436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_726
timestamp 1704896540
transform 1 0 67804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_728
timestamp 1704896540
transform 1 0 67988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_740
timestamp 1704896540
transform 1 0 69092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_752
timestamp 1704896540
transform 1 0 70196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_764
timestamp 1704896540
transform 1 0 71300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_776
timestamp 1704896540
transform 1 0 72404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_782
timestamp 1704896540
transform 1 0 72956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_784
timestamp 1704896540
transform 1 0 73140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_796
timestamp 1704896540
transform 1 0 74244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_800
timestamp 1704896540
transform 1 0 74612 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_702
timestamp 1704896540
transform 1 0 65596 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_714
timestamp 1704896540
transform 1 0 66700 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_726
timestamp 1704896540
transform 1 0 67804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_738
timestamp 1704896540
transform 1 0 68908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_750
timestamp 1704896540
transform 1 0 70012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_754
timestamp 1704896540
transform 1 0 70380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_756
timestamp 1704896540
transform 1 0 70564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_768
timestamp 1704896540
transform 1 0 71668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_780
timestamp 1704896540
transform 1 0 72772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_792
timestamp 1704896540
transform 1 0 73876 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_800
timestamp 1704896540
transform 1 0 74612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_710
timestamp 1704896540
transform 1 0 66332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_722
timestamp 1704896540
transform 1 0 67436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_726
timestamp 1704896540
transform 1 0 67804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_728
timestamp 1704896540
transform 1 0 67988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_740
timestamp 1704896540
transform 1 0 69092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_752
timestamp 1704896540
transform 1 0 70196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_764
timestamp 1704896540
transform 1 0 71300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_776
timestamp 1704896540
transform 1 0 72404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_782
timestamp 1704896540
transform 1 0 72956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_784
timestamp 1704896540
transform 1 0 73140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_796
timestamp 1704896540
transform 1 0 74244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_800
timestamp 1704896540
transform 1 0 74612 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_702
timestamp 1704896540
transform 1 0 65596 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_714
timestamp 1704896540
transform 1 0 66700 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_726
timestamp 1704896540
transform 1 0 67804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_738
timestamp 1704896540
transform 1 0 68908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_750
timestamp 1704896540
transform 1 0 70012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_754
timestamp 1704896540
transform 1 0 70380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_756
timestamp 1704896540
transform 1 0 70564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_768
timestamp 1704896540
transform 1 0 71668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_780
timestamp 1704896540
transform 1 0 72772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_792
timestamp 1704896540
transform 1 0 73876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_800
timestamp 1704896540
transform 1 0 74612 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_710
timestamp 1704896540
transform 1 0 66332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_722
timestamp 1704896540
transform 1 0 67436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_726
timestamp 1704896540
transform 1 0 67804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_728
timestamp 1704896540
transform 1 0 67988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_740
timestamp 1704896540
transform 1 0 69092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_752
timestamp 1704896540
transform 1 0 70196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_764
timestamp 1704896540
transform 1 0 71300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_776
timestamp 1704896540
transform 1 0 72404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_782
timestamp 1704896540
transform 1 0 72956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_784
timestamp 1704896540
transform 1 0 73140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_796
timestamp 1704896540
transform 1 0 74244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_800
timestamp 1704896540
transform 1 0 74612 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_702
timestamp 1704896540
transform 1 0 65596 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_714
timestamp 1704896540
transform 1 0 66700 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_726
timestamp 1704896540
transform 1 0 67804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_738
timestamp 1704896540
transform 1 0 68908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_750
timestamp 1704896540
transform 1 0 70012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_754
timestamp 1704896540
transform 1 0 70380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_756
timestamp 1704896540
transform 1 0 70564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_768
timestamp 1704896540
transform 1 0 71668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_780
timestamp 1704896540
transform 1 0 72772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_792
timestamp 1704896540
transform 1 0 73876 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_800
timestamp 1704896540
transform 1 0 74612 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_710
timestamp 1704896540
transform 1 0 66332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_722
timestamp 1704896540
transform 1 0 67436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_726
timestamp 1704896540
transform 1 0 67804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_728
timestamp 1704896540
transform 1 0 67988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_740
timestamp 1704896540
transform 1 0 69092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_752
timestamp 1704896540
transform 1 0 70196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_764
timestamp 1704896540
transform 1 0 71300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_776
timestamp 1704896540
transform 1 0 72404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_782
timestamp 1704896540
transform 1 0 72956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_784
timestamp 1704896540
transform 1 0 73140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_796
timestamp 1704896540
transform 1 0 74244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_800
timestamp 1704896540
transform 1 0 74612 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_702
timestamp 1704896540
transform 1 0 65596 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_714
timestamp 1704896540
transform 1 0 66700 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_726
timestamp 1704896540
transform 1 0 67804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_738
timestamp 1704896540
transform 1 0 68908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_750
timestamp 1704896540
transform 1 0 70012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_754
timestamp 1704896540
transform 1 0 70380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_756
timestamp 1704896540
transform 1 0 70564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_768
timestamp 1704896540
transform 1 0 71668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_780
timestamp 1704896540
transform 1 0 72772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_792
timestamp 1704896540
transform 1 0 73876 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_800
timestamp 1704896540
transform 1 0 74612 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_702
timestamp 1704896540
transform 1 0 65596 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_710
timestamp 1704896540
transform 1 0 66332 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_719
timestamp 1704896540
transform 1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_728
timestamp 1704896540
transform 1 0 67988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_740
timestamp 1704896540
transform 1 0 69092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_752
timestamp 1704896540
transform 1 0 70196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_764
timestamp 1704896540
transform 1 0 71300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_776
timestamp 1704896540
transform 1 0 72404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_782
timestamp 1704896540
transform 1 0 72956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_784
timestamp 1704896540
transform 1 0 73140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_796
timestamp 1704896540
transform 1 0 74244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_800
timestamp 1704896540
transform 1 0 74612 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_702
timestamp 1704896540
transform 1 0 65596 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_714
timestamp 1704896540
transform 1 0 66700 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_726
timestamp 1704896540
transform 1 0 67804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_738
timestamp 1704896540
transform 1 0 68908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_750
timestamp 1704896540
transform 1 0 70012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_754
timestamp 1704896540
transform 1 0 70380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_756
timestamp 1704896540
transform 1 0 70564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_768
timestamp 1704896540
transform 1 0 71668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_780
timestamp 1704896540
transform 1 0 72772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_792
timestamp 1704896540
transform 1 0 73876 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_800
timestamp 1704896540
transform 1 0 74612 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_702
timestamp 1704896540
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_714
timestamp 1704896540
transform 1 0 66700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_726
timestamp 1704896540
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_728
timestamp 1704896540
transform 1 0 67988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_740
timestamp 1704896540
transform 1 0 69092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_752
timestamp 1704896540
transform 1 0 70196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_764
timestamp 1704896540
transform 1 0 71300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_776
timestamp 1704896540
transform 1 0 72404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_782
timestamp 1704896540
transform 1 0 72956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_784
timestamp 1704896540
transform 1 0 73140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_796
timestamp 1704896540
transform 1 0 74244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_800
timestamp 1704896540
transform 1 0 74612 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_702
timestamp 1704896540
transform 1 0 65596 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_714
timestamp 1704896540
transform 1 0 66700 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_726
timestamp 1704896540
transform 1 0 67804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_738
timestamp 1704896540
transform 1 0 68908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_750
timestamp 1704896540
transform 1 0 70012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_754
timestamp 1704896540
transform 1 0 70380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_756
timestamp 1704896540
transform 1 0 70564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_768
timestamp 1704896540
transform 1 0 71668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_780
timestamp 1704896540
transform 1 0 72772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_792
timestamp 1704896540
transform 1 0 73876 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_800
timestamp 1704896540
transform 1 0 74612 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_705
timestamp 1704896540
transform 1 0 65872 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_717
timestamp 1704896540
transform 1 0 66976 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_725
timestamp 1704896540
transform 1 0 67712 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_736
timestamp 1704896540
transform 1 0 68724 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_748
timestamp 1704896540
transform 1 0 69828 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_760
timestamp 1704896540
transform 1 0 70932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_772
timestamp 1704896540
transform 1 0 72036 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_780
timestamp 1704896540
transform 1 0 72772 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_784
timestamp 1704896540
transform 1 0 73140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_796
timestamp 1704896540
transform 1 0 74244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_800
timestamp 1704896540
transform 1 0 74612 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_702
timestamp 1704896540
transform 1 0 65596 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_714
timestamp 1704896540
transform 1 0 66700 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_726
timestamp 1704896540
transform 1 0 67804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_738
timestamp 1704896540
transform 1 0 68908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_750
timestamp 1704896540
transform 1 0 70012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_754
timestamp 1704896540
transform 1 0 70380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_756
timestamp 1704896540
transform 1 0 70564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_768
timestamp 1704896540
transform 1 0 71668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_780
timestamp 1704896540
transform 1 0 72772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_792
timestamp 1704896540
transform 1 0 73876 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_800
timestamp 1704896540
transform 1 0 74612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_705
timestamp 1704896540
transform 1 0 65872 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_717
timestamp 1704896540
transform 1 0 66976 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_725
timestamp 1704896540
transform 1 0 67712 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_728
timestamp 1704896540
transform 1 0 67988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_740
timestamp 1704896540
transform 1 0 69092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_752
timestamp 1704896540
transform 1 0 70196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_764
timestamp 1704896540
transform 1 0 71300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_776
timestamp 1704896540
transform 1 0 72404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_782
timestamp 1704896540
transform 1 0 72956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_784
timestamp 1704896540
transform 1 0 73140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_796
timestamp 1704896540
transform 1 0 74244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_800
timestamp 1704896540
transform 1 0 74612 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_702
timestamp 1704896540
transform 1 0 65596 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_714
timestamp 1704896540
transform 1 0 66700 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_726
timestamp 1704896540
transform 1 0 67804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_738
timestamp 1704896540
transform 1 0 68908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_750
timestamp 1704896540
transform 1 0 70012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_754
timestamp 1704896540
transform 1 0 70380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_756
timestamp 1704896540
transform 1 0 70564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_768
timestamp 1704896540
transform 1 0 71668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_780
timestamp 1704896540
transform 1 0 72772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_792
timestamp 1704896540
transform 1 0 73876 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_800
timestamp 1704896540
transform 1 0 74612 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_702
timestamp 1704896540
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_714
timestamp 1704896540
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_726
timestamp 1704896540
transform 1 0 67804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_728
timestamp 1704896540
transform 1 0 67988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_740
timestamp 1704896540
transform 1 0 69092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_752
timestamp 1704896540
transform 1 0 70196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_764
timestamp 1704896540
transform 1 0 71300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_776
timestamp 1704896540
transform 1 0 72404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_782
timestamp 1704896540
transform 1 0 72956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_784
timestamp 1704896540
transform 1 0 73140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_796
timestamp 1704896540
transform 1 0 74244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_800
timestamp 1704896540
transform 1 0 74612 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_702
timestamp 1704896540
transform 1 0 65596 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_714
timestamp 1704896540
transform 1 0 66700 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_726
timestamp 1704896540
transform 1 0 67804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_738
timestamp 1704896540
transform 1 0 68908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_750
timestamp 1704896540
transform 1 0 70012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_754
timestamp 1704896540
transform 1 0 70380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_756
timestamp 1704896540
transform 1 0 70564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_768
timestamp 1704896540
transform 1 0 71668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_780
timestamp 1704896540
transform 1 0 72772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_792
timestamp 1704896540
transform 1 0 73876 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_800
timestamp 1704896540
transform 1 0 74612 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_702
timestamp 1704896540
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_714
timestamp 1704896540
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_726
timestamp 1704896540
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_728
timestamp 1704896540
transform 1 0 67988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_740
timestamp 1704896540
transform 1 0 69092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_752
timestamp 1704896540
transform 1 0 70196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_764
timestamp 1704896540
transform 1 0 71300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_776
timestamp 1704896540
transform 1 0 72404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_782
timestamp 1704896540
transform 1 0 72956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_784
timestamp 1704896540
transform 1 0 73140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_796
timestamp 1704896540
transform 1 0 74244 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_800
timestamp 1704896540
transform 1 0 74612 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_702
timestamp 1704896540
transform 1 0 65596 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_714
timestamp 1704896540
transform 1 0 66700 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_726
timestamp 1704896540
transform 1 0 67804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_738
timestamp 1704896540
transform 1 0 68908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_750
timestamp 1704896540
transform 1 0 70012 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_754
timestamp 1704896540
transform 1 0 70380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_756
timestamp 1704896540
transform 1 0 70564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_768
timestamp 1704896540
transform 1 0 71668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_780
timestamp 1704896540
transform 1 0 72772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_792
timestamp 1704896540
transform 1 0 73876 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_800
timestamp 1704896540
transform 1 0 74612 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_708
timestamp 1704896540
transform 1 0 66148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_720
timestamp 1704896540
transform 1 0 67252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_726
timestamp 1704896540
transform 1 0 67804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_728
timestamp 1704896540
transform 1 0 67988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_740
timestamp 1704896540
transform 1 0 69092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_752
timestamp 1704896540
transform 1 0 70196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_764
timestamp 1704896540
transform 1 0 71300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_776
timestamp 1704896540
transform 1 0 72404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_782
timestamp 1704896540
transform 1 0 72956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_784
timestamp 1704896540
transform 1 0 73140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_84_796
timestamp 1704896540
transform 1 0 74244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_800
timestamp 1704896540
transform 1 0 74612 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_702
timestamp 1704896540
transform 1 0 65596 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_714
timestamp 1704896540
transform 1 0 66700 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_726
timestamp 1704896540
transform 1 0 67804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_738
timestamp 1704896540
transform 1 0 68908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_750
timestamp 1704896540
transform 1 0 70012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_754
timestamp 1704896540
transform 1 0 70380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_756
timestamp 1704896540
transform 1 0 70564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_768
timestamp 1704896540
transform 1 0 71668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_780
timestamp 1704896540
transform 1 0 72772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_792
timestamp 1704896540
transform 1 0 73876 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_800
timestamp 1704896540
transform 1 0 74612 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_702
timestamp 1704896540
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_714
timestamp 1704896540
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_726
timestamp 1704896540
transform 1 0 67804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_728
timestamp 1704896540
transform 1 0 67988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_740
timestamp 1704896540
transform 1 0 69092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_752
timestamp 1704896540
transform 1 0 70196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_764
timestamp 1704896540
transform 1 0 71300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_776
timestamp 1704896540
transform 1 0 72404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_782
timestamp 1704896540
transform 1 0 72956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_784
timestamp 1704896540
transform 1 0 73140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86_796
timestamp 1704896540
transform 1 0 74244 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_800
timestamp 1704896540
transform 1 0 74612 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_702
timestamp 1704896540
transform 1 0 65596 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_714
timestamp 1704896540
transform 1 0 66700 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_726
timestamp 1704896540
transform 1 0 67804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_738
timestamp 1704896540
transform 1 0 68908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_750
timestamp 1704896540
transform 1 0 70012 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_754
timestamp 1704896540
transform 1 0 70380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_756
timestamp 1704896540
transform 1 0 70564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_768
timestamp 1704896540
transform 1 0 71668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_780
timestamp 1704896540
transform 1 0 72772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_792
timestamp 1704896540
transform 1 0 73876 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_800
timestamp 1704896540
transform 1 0 74612 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_705
timestamp 1704896540
transform 1 0 65872 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_717
timestamp 1704896540
transform 1 0 66976 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88_725
timestamp 1704896540
transform 1 0 67712 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_728
timestamp 1704896540
transform 1 0 67988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_740
timestamp 1704896540
transform 1 0 69092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_752
timestamp 1704896540
transform 1 0 70196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_764
timestamp 1704896540
transform 1 0 71300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_776
timestamp 1704896540
transform 1 0 72404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_782
timestamp 1704896540
transform 1 0 72956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_784
timestamp 1704896540
transform 1 0 73140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88_796
timestamp 1704896540
transform 1 0 74244 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_800
timestamp 1704896540
transform 1 0 74612 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_705
timestamp 1704896540
transform 1 0 65872 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_717
timestamp 1704896540
transform 1 0 66976 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_729
timestamp 1704896540
transform 1 0 68080 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_741
timestamp 1704896540
transform 1 0 69184 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_753
timestamp 1704896540
transform 1 0 70288 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_756
timestamp 1704896540
transform 1 0 70564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_768
timestamp 1704896540
transform 1 0 71668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_780
timestamp 1704896540
transform 1 0 72772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_792
timestamp 1704896540
transform 1 0 73876 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_800
timestamp 1704896540
transform 1 0 74612 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_705
timestamp 1704896540
transform 1 0 65872 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_717
timestamp 1704896540
transform 1 0 66976 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_725
timestamp 1704896540
transform 1 0 67712 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_728
timestamp 1704896540
transform 1 0 67988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_740
timestamp 1704896540
transform 1 0 69092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_752
timestamp 1704896540
transform 1 0 70196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_764
timestamp 1704896540
transform 1 0 71300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_776
timestamp 1704896540
transform 1 0 72404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_782
timestamp 1704896540
transform 1 0 72956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_784
timestamp 1704896540
transform 1 0 73140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90_796
timestamp 1704896540
transform 1 0 74244 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_800
timestamp 1704896540
transform 1 0 74612 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_702
timestamp 1704896540
transform 1 0 65596 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_714
timestamp 1704896540
transform 1 0 66700 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_726
timestamp 1704896540
transform 1 0 67804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_738
timestamp 1704896540
transform 1 0 68908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_750
timestamp 1704896540
transform 1 0 70012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_754
timestamp 1704896540
transform 1 0 70380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_756
timestamp 1704896540
transform 1 0 70564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_768
timestamp 1704896540
transform 1 0 71668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_780
timestamp 1704896540
transform 1 0 72772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_792
timestamp 1704896540
transform 1 0 73876 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_800
timestamp 1704896540
transform 1 0 74612 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_702
timestamp 1704896540
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_714
timestamp 1704896540
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_726
timestamp 1704896540
transform 1 0 67804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_728
timestamp 1704896540
transform 1 0 67988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_740
timestamp 1704896540
transform 1 0 69092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_752
timestamp 1704896540
transform 1 0 70196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_764
timestamp 1704896540
transform 1 0 71300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_776
timestamp 1704896540
transform 1 0 72404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_782
timestamp 1704896540
transform 1 0 72956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_784
timestamp 1704896540
transform 1 0 73140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92_796
timestamp 1704896540
transform 1 0 74244 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_800
timestamp 1704896540
transform 1 0 74612 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_702
timestamp 1704896540
transform 1 0 65596 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_714
timestamp 1704896540
transform 1 0 66700 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_726
timestamp 1704896540
transform 1 0 67804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_738
timestamp 1704896540
transform 1 0 68908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_750
timestamp 1704896540
transform 1 0 70012 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_754
timestamp 1704896540
transform 1 0 70380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_756
timestamp 1704896540
transform 1 0 70564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_768
timestamp 1704896540
transform 1 0 71668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_780
timestamp 1704896540
transform 1 0 72772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_792
timestamp 1704896540
transform 1 0 73876 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_800
timestamp 1704896540
transform 1 0 74612 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_708
timestamp 1704896540
transform 1 0 66148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_720
timestamp 1704896540
transform 1 0 67252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_726
timestamp 1704896540
transform 1 0 67804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_728
timestamp 1704896540
transform 1 0 67988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_740
timestamp 1704896540
transform 1 0 69092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_752
timestamp 1704896540
transform 1 0 70196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_764
timestamp 1704896540
transform 1 0 71300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_776
timestamp 1704896540
transform 1 0 72404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_782
timestamp 1704896540
transform 1 0 72956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_784
timestamp 1704896540
transform 1 0 73140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_796
timestamp 1704896540
transform 1 0 74244 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_800
timestamp 1704896540
transform 1 0 74612 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_702
timestamp 1704896540
transform 1 0 65596 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_714
timestamp 1704896540
transform 1 0 66700 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_726
timestamp 1704896540
transform 1 0 67804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_738
timestamp 1704896540
transform 1 0 68908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_750
timestamp 1704896540
transform 1 0 70012 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_754
timestamp 1704896540
transform 1 0 70380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_756
timestamp 1704896540
transform 1 0 70564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_768
timestamp 1704896540
transform 1 0 71668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_780
timestamp 1704896540
transform 1 0 72772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_792
timestamp 1704896540
transform 1 0 73876 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_800
timestamp 1704896540
transform 1 0 74612 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_702
timestamp 1704896540
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_714
timestamp 1704896540
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_726
timestamp 1704896540
transform 1 0 67804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_728
timestamp 1704896540
transform 1 0 67988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_740
timestamp 1704896540
transform 1 0 69092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_752
timestamp 1704896540
transform 1 0 70196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_764
timestamp 1704896540
transform 1 0 71300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_776
timestamp 1704896540
transform 1 0 72404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_782
timestamp 1704896540
transform 1 0 72956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_784
timestamp 1704896540
transform 1 0 73140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_796
timestamp 1704896540
transform 1 0 74244 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_800
timestamp 1704896540
transform 1 0 74612 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_702
timestamp 1704896540
transform 1 0 65596 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_714
timestamp 1704896540
transform 1 0 66700 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_726
timestamp 1704896540
transform 1 0 67804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_738
timestamp 1704896540
transform 1 0 68908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_750
timestamp 1704896540
transform 1 0 70012 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_754
timestamp 1704896540
transform 1 0 70380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_756
timestamp 1704896540
transform 1 0 70564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_768
timestamp 1704896540
transform 1 0 71668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_780
timestamp 1704896540
transform 1 0 72772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_792
timestamp 1704896540
transform 1 0 73876 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_800
timestamp 1704896540
transform 1 0 74612 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_702
timestamp 1704896540
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_714
timestamp 1704896540
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_726
timestamp 1704896540
transform 1 0 67804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_728
timestamp 1704896540
transform 1 0 67988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_740
timestamp 1704896540
transform 1 0 69092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_752
timestamp 1704896540
transform 1 0 70196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_764
timestamp 1704896540
transform 1 0 71300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_776
timestamp 1704896540
transform 1 0 72404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_782
timestamp 1704896540
transform 1 0 72956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_784
timestamp 1704896540
transform 1 0 73140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_796
timestamp 1704896540
transform 1 0 74244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_800
timestamp 1704896540
transform 1 0 74612 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_702
timestamp 1704896540
transform 1 0 65596 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_714
timestamp 1704896540
transform 1 0 66700 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_726
timestamp 1704896540
transform 1 0 67804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_738
timestamp 1704896540
transform 1 0 68908 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_750
timestamp 1704896540
transform 1 0 70012 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_754
timestamp 1704896540
transform 1 0 70380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_756
timestamp 1704896540
transform 1 0 70564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_768
timestamp 1704896540
transform 1 0 71668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_780
timestamp 1704896540
transform 1 0 72772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_792
timestamp 1704896540
transform 1 0 73876 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_800
timestamp 1704896540
transform 1 0 74612 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_702
timestamp 1704896540
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_714
timestamp 1704896540
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_726
timestamp 1704896540
transform 1 0 67804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_728
timestamp 1704896540
transform 1 0 67988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_740
timestamp 1704896540
transform 1 0 69092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_752
timestamp 1704896540
transform 1 0 70196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_764
timestamp 1704896540
transform 1 0 71300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_776
timestamp 1704896540
transform 1 0 72404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_782
timestamp 1704896540
transform 1 0 72956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_784
timestamp 1704896540
transform 1 0 73140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_796
timestamp 1704896540
transform 1 0 74244 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_800
timestamp 1704896540
transform 1 0 74612 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_702
timestamp 1704896540
transform 1 0 65596 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_714
timestamp 1704896540
transform 1 0 66700 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_726
timestamp 1704896540
transform 1 0 67804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_738
timestamp 1704896540
transform 1 0 68908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_750
timestamp 1704896540
transform 1 0 70012 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_754
timestamp 1704896540
transform 1 0 70380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_756
timestamp 1704896540
transform 1 0 70564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_768
timestamp 1704896540
transform 1 0 71668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_780
timestamp 1704896540
transform 1 0 72772 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_792
timestamp 1704896540
transform 1 0 73876 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_800
timestamp 1704896540
transform 1 0 74612 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_702
timestamp 1704896540
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_714
timestamp 1704896540
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_726
timestamp 1704896540
transform 1 0 67804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_728
timestamp 1704896540
transform 1 0 67988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_740
timestamp 1704896540
transform 1 0 69092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_752
timestamp 1704896540
transform 1 0 70196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_764
timestamp 1704896540
transform 1 0 71300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_776
timestamp 1704896540
transform 1 0 72404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_782
timestamp 1704896540
transform 1 0 72956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_784
timestamp 1704896540
transform 1 0 73140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_796
timestamp 1704896540
transform 1 0 74244 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_800
timestamp 1704896540
transform 1 0 74612 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_702
timestamp 1704896540
transform 1 0 65596 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_714
timestamp 1704896540
transform 1 0 66700 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_726
timestamp 1704896540
transform 1 0 67804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_738
timestamp 1704896540
transform 1 0 68908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_750
timestamp 1704896540
transform 1 0 70012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_754
timestamp 1704896540
transform 1 0 70380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_756
timestamp 1704896540
transform 1 0 70564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_768
timestamp 1704896540
transform 1 0 71668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_780
timestamp 1704896540
transform 1 0 72772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_792
timestamp 1704896540
transform 1 0 73876 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_800
timestamp 1704896540
transform 1 0 74612 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_702
timestamp 1704896540
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_714
timestamp 1704896540
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_726
timestamp 1704896540
transform 1 0 67804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_728
timestamp 1704896540
transform 1 0 67988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_740
timestamp 1704896540
transform 1 0 69092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_752
timestamp 1704896540
transform 1 0 70196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_764
timestamp 1704896540
transform 1 0 71300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_776
timestamp 1704896540
transform 1 0 72404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_782
timestamp 1704896540
transform 1 0 72956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_784
timestamp 1704896540
transform 1 0 73140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_796
timestamp 1704896540
transform 1 0 74244 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_800
timestamp 1704896540
transform 1 0 74612 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_702
timestamp 1704896540
transform 1 0 65596 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_714
timestamp 1704896540
transform 1 0 66700 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_726
timestamp 1704896540
transform 1 0 67804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_738
timestamp 1704896540
transform 1 0 68908 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_750
timestamp 1704896540
transform 1 0 70012 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_754
timestamp 1704896540
transform 1 0 70380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_756
timestamp 1704896540
transform 1 0 70564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_768
timestamp 1704896540
transform 1 0 71668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_780
timestamp 1704896540
transform 1 0 72772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_792
timestamp 1704896540
transform 1 0 73876 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_800
timestamp 1704896540
transform 1 0 74612 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_702
timestamp 1704896540
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_714
timestamp 1704896540
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_726
timestamp 1704896540
transform 1 0 67804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_728
timestamp 1704896540
transform 1 0 67988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_740
timestamp 1704896540
transform 1 0 69092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_752
timestamp 1704896540
transform 1 0 70196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_764
timestamp 1704896540
transform 1 0 71300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_776
timestamp 1704896540
transform 1 0 72404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_782
timestamp 1704896540
transform 1 0 72956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_784
timestamp 1704896540
transform 1 0 73140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106_796
timestamp 1704896540
transform 1 0 74244 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_800
timestamp 1704896540
transform 1 0 74612 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_702
timestamp 1704896540
transform 1 0 65596 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_714
timestamp 1704896540
transform 1 0 66700 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_726
timestamp 1704896540
transform 1 0 67804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_738
timestamp 1704896540
transform 1 0 68908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_750
timestamp 1704896540
transform 1 0 70012 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_754
timestamp 1704896540
transform 1 0 70380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_756
timestamp 1704896540
transform 1 0 70564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_768
timestamp 1704896540
transform 1 0 71668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_780
timestamp 1704896540
transform 1 0 72772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_792
timestamp 1704896540
transform 1 0 73876 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_800
timestamp 1704896540
transform 1 0 74612 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_702
timestamp 1704896540
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_714
timestamp 1704896540
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_726
timestamp 1704896540
transform 1 0 67804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_728
timestamp 1704896540
transform 1 0 67988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_740
timestamp 1704896540
transform 1 0 69092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_752
timestamp 1704896540
transform 1 0 70196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_764
timestamp 1704896540
transform 1 0 71300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_776
timestamp 1704896540
transform 1 0 72404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_782
timestamp 1704896540
transform 1 0 72956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_784
timestamp 1704896540
transform 1 0 73140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108_796
timestamp 1704896540
transform 1 0 74244 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_800
timestamp 1704896540
transform 1 0 74612 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_702
timestamp 1704896540
transform 1 0 65596 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_714
timestamp 1704896540
transform 1 0 66700 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_726
timestamp 1704896540
transform 1 0 67804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_738
timestamp 1704896540
transform 1 0 68908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_750
timestamp 1704896540
transform 1 0 70012 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_754
timestamp 1704896540
transform 1 0 70380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_756
timestamp 1704896540
transform 1 0 70564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_768
timestamp 1704896540
transform 1 0 71668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_780
timestamp 1704896540
transform 1 0 72772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_792
timestamp 1704896540
transform 1 0 73876 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_800
timestamp 1704896540
transform 1 0 74612 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_702
timestamp 1704896540
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_714
timestamp 1704896540
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_726
timestamp 1704896540
transform 1 0 67804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_728
timestamp 1704896540
transform 1 0 67988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_740
timestamp 1704896540
transform 1 0 69092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_752
timestamp 1704896540
transform 1 0 70196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_764
timestamp 1704896540
transform 1 0 71300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_776
timestamp 1704896540
transform 1 0 72404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_782
timestamp 1704896540
transform 1 0 72956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_784
timestamp 1704896540
transform 1 0 73140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_796
timestamp 1704896540
transform 1 0 74244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_800
timestamp 1704896540
transform 1 0 74612 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_702
timestamp 1704896540
transform 1 0 65596 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_714
timestamp 1704896540
transform 1 0 66700 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_726
timestamp 1704896540
transform 1 0 67804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_738
timestamp 1704896540
transform 1 0 68908 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_750
timestamp 1704896540
transform 1 0 70012 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_754
timestamp 1704896540
transform 1 0 70380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_756
timestamp 1704896540
transform 1 0 70564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_768
timestamp 1704896540
transform 1 0 71668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_780
timestamp 1704896540
transform 1 0 72772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_792
timestamp 1704896540
transform 1 0 73876 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_800
timestamp 1704896540
transform 1 0 74612 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_702
timestamp 1704896540
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_714
timestamp 1704896540
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_726
timestamp 1704896540
transform 1 0 67804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_728
timestamp 1704896540
transform 1 0 67988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_740
timestamp 1704896540
transform 1 0 69092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_752
timestamp 1704896540
transform 1 0 70196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_764
timestamp 1704896540
transform 1 0 71300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_776
timestamp 1704896540
transform 1 0 72404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_782
timestamp 1704896540
transform 1 0 72956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_784
timestamp 1704896540
transform 1 0 73140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_796
timestamp 1704896540
transform 1 0 74244 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_800
timestamp 1704896540
transform 1 0 74612 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_702
timestamp 1704896540
transform 1 0 65596 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_714
timestamp 1704896540
transform 1 0 66700 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_726
timestamp 1704896540
transform 1 0 67804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_738
timestamp 1704896540
transform 1 0 68908 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_750
timestamp 1704896540
transform 1 0 70012 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_754
timestamp 1704896540
transform 1 0 70380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_756
timestamp 1704896540
transform 1 0 70564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_768
timestamp 1704896540
transform 1 0 71668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_780
timestamp 1704896540
transform 1 0 72772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_792
timestamp 1704896540
transform 1 0 73876 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_800
timestamp 1704896540
transform 1 0 74612 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_702
timestamp 1704896540
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_714
timestamp 1704896540
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_726
timestamp 1704896540
transform 1 0 67804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_728
timestamp 1704896540
transform 1 0 67988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_740
timestamp 1704896540
transform 1 0 69092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_752
timestamp 1704896540
transform 1 0 70196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_764
timestamp 1704896540
transform 1 0 71300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_776
timestamp 1704896540
transform 1 0 72404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_782
timestamp 1704896540
transform 1 0 72956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_784
timestamp 1704896540
transform 1 0 73140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_796
timestamp 1704896540
transform 1 0 74244 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_800
timestamp 1704896540
transform 1 0 74612 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_702
timestamp 1704896540
transform 1 0 65596 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_714
timestamp 1704896540
transform 1 0 66700 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_726
timestamp 1704896540
transform 1 0 67804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_738
timestamp 1704896540
transform 1 0 68908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_750
timestamp 1704896540
transform 1 0 70012 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_754
timestamp 1704896540
transform 1 0 70380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_756
timestamp 1704896540
transform 1 0 70564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_768
timestamp 1704896540
transform 1 0 71668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_780
timestamp 1704896540
transform 1 0 72772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_792
timestamp 1704896540
transform 1 0 73876 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_800
timestamp 1704896540
transform 1 0 74612 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_702
timestamp 1704896540
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_714
timestamp 1704896540
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_726
timestamp 1704896540
transform 1 0 67804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_728
timestamp 1704896540
transform 1 0 67988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_740
timestamp 1704896540
transform 1 0 69092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_752
timestamp 1704896540
transform 1 0 70196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_764
timestamp 1704896540
transform 1 0 71300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_776
timestamp 1704896540
transform 1 0 72404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_782
timestamp 1704896540
transform 1 0 72956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_784
timestamp 1704896540
transform 1 0 73140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_796
timestamp 1704896540
transform 1 0 74244 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_800
timestamp 1704896540
transform 1 0 74612 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_702
timestamp 1704896540
transform 1 0 65596 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_714
timestamp 1704896540
transform 1 0 66700 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_726
timestamp 1704896540
transform 1 0 67804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_738
timestamp 1704896540
transform 1 0 68908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_750
timestamp 1704896540
transform 1 0 70012 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_754
timestamp 1704896540
transform 1 0 70380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_756
timestamp 1704896540
transform 1 0 70564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_768
timestamp 1704896540
transform 1 0 71668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_780
timestamp 1704896540
transform 1 0 72772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_792
timestamp 1704896540
transform 1 0 73876 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_800
timestamp 1704896540
transform 1 0 74612 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_702
timestamp 1704896540
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_714
timestamp 1704896540
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_726
timestamp 1704896540
transform 1 0 67804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_728
timestamp 1704896540
transform 1 0 67988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_740
timestamp 1704896540
transform 1 0 69092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_752
timestamp 1704896540
transform 1 0 70196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_764
timestamp 1704896540
transform 1 0 71300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_776
timestamp 1704896540
transform 1 0 72404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_782
timestamp 1704896540
transform 1 0 72956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_784
timestamp 1704896540
transform 1 0 73140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_796
timestamp 1704896540
transform 1 0 74244 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_800
timestamp 1704896540
transform 1 0 74612 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_702
timestamp 1704896540
transform 1 0 65596 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_714
timestamp 1704896540
transform 1 0 66700 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_726
timestamp 1704896540
transform 1 0 67804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_738
timestamp 1704896540
transform 1 0 68908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_750
timestamp 1704896540
transform 1 0 70012 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_754
timestamp 1704896540
transform 1 0 70380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_756
timestamp 1704896540
transform 1 0 70564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_768
timestamp 1704896540
transform 1 0 71668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_780
timestamp 1704896540
transform 1 0 72772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_792
timestamp 1704896540
transform 1 0 73876 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_800
timestamp 1704896540
transform 1 0 74612 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_702
timestamp 1704896540
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_714
timestamp 1704896540
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_726
timestamp 1704896540
transform 1 0 67804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_728
timestamp 1704896540
transform 1 0 67988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_740
timestamp 1704896540
transform 1 0 69092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_752
timestamp 1704896540
transform 1 0 70196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_764
timestamp 1704896540
transform 1 0 71300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_776
timestamp 1704896540
transform 1 0 72404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_782
timestamp 1704896540
transform 1 0 72956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_784
timestamp 1704896540
transform 1 0 73140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_796
timestamp 1704896540
transform 1 0 74244 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_800
timestamp 1704896540
transform 1 0 74612 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_702
timestamp 1704896540
transform 1 0 65596 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_714
timestamp 1704896540
transform 1 0 66700 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_726
timestamp 1704896540
transform 1 0 67804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_738
timestamp 1704896540
transform 1 0 68908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_750
timestamp 1704896540
transform 1 0 70012 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_754
timestamp 1704896540
transform 1 0 70380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_756
timestamp 1704896540
transform 1 0 70564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_768
timestamp 1704896540
transform 1 0 71668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_780
timestamp 1704896540
transform 1 0 72772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_792
timestamp 1704896540
transform 1 0 73876 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_800
timestamp 1704896540
transform 1 0 74612 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_702
timestamp 1704896540
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_714
timestamp 1704896540
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_726
timestamp 1704896540
transform 1 0 67804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_728
timestamp 1704896540
transform 1 0 67988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_740
timestamp 1704896540
transform 1 0 69092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_752
timestamp 1704896540
transform 1 0 70196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_764
timestamp 1704896540
transform 1 0 71300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_776
timestamp 1704896540
transform 1 0 72404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_782
timestamp 1704896540
transform 1 0 72956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_784
timestamp 1704896540
transform 1 0 73140 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_796
timestamp 1704896540
transform 1 0 74244 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_800
timestamp 1704896540
transform 1 0 74612 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_702
timestamp 1704896540
transform 1 0 65596 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_714
timestamp 1704896540
transform 1 0 66700 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_726
timestamp 1704896540
transform 1 0 67804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_738
timestamp 1704896540
transform 1 0 68908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_750
timestamp 1704896540
transform 1 0 70012 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_754
timestamp 1704896540
transform 1 0 70380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_756
timestamp 1704896540
transform 1 0 70564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_768
timestamp 1704896540
transform 1 0 71668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_780
timestamp 1704896540
transform 1 0 72772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_792
timestamp 1704896540
transform 1 0 73876 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_800
timestamp 1704896540
transform 1 0 74612 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_702
timestamp 1704896540
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_714
timestamp 1704896540
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_726
timestamp 1704896540
transform 1 0 67804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_728
timestamp 1704896540
transform 1 0 67988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_740
timestamp 1704896540
transform 1 0 69092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_752
timestamp 1704896540
transform 1 0 70196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_764
timestamp 1704896540
transform 1 0 71300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_124_776
timestamp 1704896540
transform 1 0 72404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_782
timestamp 1704896540
transform 1 0 72956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_784
timestamp 1704896540
transform 1 0 73140 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124_796
timestamp 1704896540
transform 1 0 74244 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_800
timestamp 1704896540
transform 1 0 74612 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_702
timestamp 1704896540
transform 1 0 65596 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_714
timestamp 1704896540
transform 1 0 66700 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_726
timestamp 1704896540
transform 1 0 67804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_738
timestamp 1704896540
transform 1 0 68908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125_750
timestamp 1704896540
transform 1 0 70012 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_754
timestamp 1704896540
transform 1 0 70380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_756
timestamp 1704896540
transform 1 0 70564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_768
timestamp 1704896540
transform 1 0 71668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_780
timestamp 1704896540
transform 1 0 72772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_792
timestamp 1704896540
transform 1 0 73876 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_800
timestamp 1704896540
transform 1 0 74612 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_702
timestamp 1704896540
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_714
timestamp 1704896540
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_726
timestamp 1704896540
transform 1 0 67804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_728
timestamp 1704896540
transform 1 0 67988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_740
timestamp 1704896540
transform 1 0 69092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_752
timestamp 1704896540
transform 1 0 70196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_764
timestamp 1704896540
transform 1 0 71300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_126_776
timestamp 1704896540
transform 1 0 72404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_782
timestamp 1704896540
transform 1 0 72956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_784
timestamp 1704896540
transform 1 0 73140 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126_796
timestamp 1704896540
transform 1 0 74244 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_800
timestamp 1704896540
transform 1 0 74612 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_702
timestamp 1704896540
transform 1 0 65596 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_714
timestamp 1704896540
transform 1 0 66700 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_726
timestamp 1704896540
transform 1 0 67804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_738
timestamp 1704896540
transform 1 0 68908 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127_750
timestamp 1704896540
transform 1 0 70012 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_754
timestamp 1704896540
transform 1 0 70380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_756
timestamp 1704896540
transform 1 0 70564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_768
timestamp 1704896540
transform 1 0 71668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_780
timestamp 1704896540
transform 1 0 72772 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_792
timestamp 1704896540
transform 1 0 73876 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_800
timestamp 1704896540
transform 1 0 74612 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_702
timestamp 1704896540
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_714
timestamp 1704896540
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_726
timestamp 1704896540
transform 1 0 67804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_728
timestamp 1704896540
transform 1 0 67988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_740
timestamp 1704896540
transform 1 0 69092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_752
timestamp 1704896540
transform 1 0 70196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_764
timestamp 1704896540
transform 1 0 71300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_128_776
timestamp 1704896540
transform 1 0 72404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_782
timestamp 1704896540
transform 1 0 72956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_784
timestamp 1704896540
transform 1 0 73140 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128_796
timestamp 1704896540
transform 1 0 74244 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_800
timestamp 1704896540
transform 1 0 74612 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_702
timestamp 1704896540
transform 1 0 65596 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_714
timestamp 1704896540
transform 1 0 66700 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_726
timestamp 1704896540
transform 1 0 67804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_738
timestamp 1704896540
transform 1 0 68908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129_750
timestamp 1704896540
transform 1 0 70012 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_754
timestamp 1704896540
transform 1 0 70380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_756
timestamp 1704896540
transform 1 0 70564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_768
timestamp 1704896540
transform 1 0 71668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_780
timestamp 1704896540
transform 1 0 72772 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_792
timestamp 1704896540
transform 1 0 73876 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_800
timestamp 1704896540
transform 1 0 74612 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_702
timestamp 1704896540
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_714
timestamp 1704896540
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_726
timestamp 1704896540
transform 1 0 67804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_728
timestamp 1704896540
transform 1 0 67988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_740
timestamp 1704896540
transform 1 0 69092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_752
timestamp 1704896540
transform 1 0 70196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_764
timestamp 1704896540
transform 1 0 71300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_130_776
timestamp 1704896540
transform 1 0 72404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_782
timestamp 1704896540
transform 1 0 72956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_784
timestamp 1704896540
transform 1 0 73140 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130_796
timestamp 1704896540
transform 1 0 74244 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_800
timestamp 1704896540
transform 1 0 74612 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_702
timestamp 1704896540
transform 1 0 65596 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_714
timestamp 1704896540
transform 1 0 66700 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_726
timestamp 1704896540
transform 1 0 67804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_738
timestamp 1704896540
transform 1 0 68908 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131_750
timestamp 1704896540
transform 1 0 70012 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_754
timestamp 1704896540
transform 1 0 70380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_756
timestamp 1704896540
transform 1 0 70564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_768
timestamp 1704896540
transform 1 0 71668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_780
timestamp 1704896540
transform 1 0 72772 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_792
timestamp 1704896540
transform 1 0 73876 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_800
timestamp 1704896540
transform 1 0 74612 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_702
timestamp 1704896540
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_714
timestamp 1704896540
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_726
timestamp 1704896540
transform 1 0 67804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_728
timestamp 1704896540
transform 1 0 67988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_740
timestamp 1704896540
transform 1 0 69092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_752
timestamp 1704896540
transform 1 0 70196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_764
timestamp 1704896540
transform 1 0 71300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_132_776
timestamp 1704896540
transform 1 0 72404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_782
timestamp 1704896540
transform 1 0 72956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_784
timestamp 1704896540
transform 1 0 73140 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132_796
timestamp 1704896540
transform 1 0 74244 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_800
timestamp 1704896540
transform 1 0 74612 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_702
timestamp 1704896540
transform 1 0 65596 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_714
timestamp 1704896540
transform 1 0 66700 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_726
timestamp 1704896540
transform 1 0 67804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_738
timestamp 1704896540
transform 1 0 68908 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_750
timestamp 1704896540
transform 1 0 70012 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_754
timestamp 1704896540
transform 1 0 70380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_756
timestamp 1704896540
transform 1 0 70564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_768
timestamp 1704896540
transform 1 0 71668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_780
timestamp 1704896540
transform 1 0 72772 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_792
timestamp 1704896540
transform 1 0 73876 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_800
timestamp 1704896540
transform 1 0 74612 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_702
timestamp 1704896540
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_714
timestamp 1704896540
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_726
timestamp 1704896540
transform 1 0 67804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_728
timestamp 1704896540
transform 1 0 67988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_740
timestamp 1704896540
transform 1 0 69092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_752
timestamp 1704896540
transform 1 0 70196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_764
timestamp 1704896540
transform 1 0 71300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134_776
timestamp 1704896540
transform 1 0 72404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_782
timestamp 1704896540
transform 1 0 72956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_784
timestamp 1704896540
transform 1 0 73140 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134_796
timestamp 1704896540
transform 1 0 74244 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_800
timestamp 1704896540
transform 1 0 74612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_702
timestamp 1704896540
transform 1 0 65596 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_714
timestamp 1704896540
transform 1 0 66700 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_726
timestamp 1704896540
transform 1 0 67804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_738
timestamp 1704896540
transform 1 0 68908 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135_750
timestamp 1704896540
transform 1 0 70012 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_754
timestamp 1704896540
transform 1 0 70380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_756
timestamp 1704896540
transform 1 0 70564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_768
timestamp 1704896540
transform 1 0 71668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_780
timestamp 1704896540
transform 1 0 72772 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_792
timestamp 1704896540
transform 1 0 73876 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_800
timestamp 1704896540
transform 1 0 74612 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_702
timestamp 1704896540
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_714
timestamp 1704896540
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_726
timestamp 1704896540
transform 1 0 67804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_728
timestamp 1704896540
transform 1 0 67988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_740
timestamp 1704896540
transform 1 0 69092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_752
timestamp 1704896540
transform 1 0 70196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_764
timestamp 1704896540
transform 1 0 71300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_136_776
timestamp 1704896540
transform 1 0 72404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_782
timestamp 1704896540
transform 1 0 72956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_784
timestamp 1704896540
transform 1 0 73140 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136_796
timestamp 1704896540
transform 1 0 74244 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_800
timestamp 1704896540
transform 1 0 74612 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_702
timestamp 1704896540
transform 1 0 65596 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_714
timestamp 1704896540
transform 1 0 66700 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_726
timestamp 1704896540
transform 1 0 67804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_738
timestamp 1704896540
transform 1 0 68908 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137_750
timestamp 1704896540
transform 1 0 70012 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_754
timestamp 1704896540
transform 1 0 70380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_756
timestamp 1704896540
transform 1 0 70564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_768
timestamp 1704896540
transform 1 0 71668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_780
timestamp 1704896540
transform 1 0 72772 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_792
timestamp 1704896540
transform 1 0 73876 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_800
timestamp 1704896540
transform 1 0 74612 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_702
timestamp 1704896540
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_714
timestamp 1704896540
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_726
timestamp 1704896540
transform 1 0 67804 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_728
timestamp 1704896540
transform 1 0 67988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_740
timestamp 1704896540
transform 1 0 69092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_752
timestamp 1704896540
transform 1 0 70196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_764
timestamp 1704896540
transform 1 0 71300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_138_776
timestamp 1704896540
transform 1 0 72404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_782
timestamp 1704896540
transform 1 0 72956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_784
timestamp 1704896540
transform 1 0 73140 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_138_796
timestamp 1704896540
transform 1 0 74244 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_800
timestamp 1704896540
transform 1 0 74612 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_702
timestamp 1704896540
transform 1 0 65596 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_714
timestamp 1704896540
transform 1 0 66700 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_726
timestamp 1704896540
transform 1 0 67804 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_738
timestamp 1704896540
transform 1 0 68908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_139_750
timestamp 1704896540
transform 1 0 70012 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_754
timestamp 1704896540
transform 1 0 70380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_756
timestamp 1704896540
transform 1 0 70564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_768
timestamp 1704896540
transform 1 0 71668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_780
timestamp 1704896540
transform 1 0 72772 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_139_792
timestamp 1704896540
transform 1 0 73876 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_800
timestamp 1704896540
transform 1 0 74612 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_702
timestamp 1704896540
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_714
timestamp 1704896540
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_726
timestamp 1704896540
transform 1 0 67804 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_728
timestamp 1704896540
transform 1 0 67988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_740
timestamp 1704896540
transform 1 0 69092 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_752
timestamp 1704896540
transform 1 0 70196 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_764
timestamp 1704896540
transform 1 0 71300 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_140_776
timestamp 1704896540
transform 1 0 72404 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_782
timestamp 1704896540
transform 1 0 72956 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_784
timestamp 1704896540
transform 1 0 73140 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140_796
timestamp 1704896540
transform 1 0 74244 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_800
timestamp 1704896540
transform 1 0 74612 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_702
timestamp 1704896540
transform 1 0 65596 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_714
timestamp 1704896540
transform 1 0 66700 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_726
timestamp 1704896540
transform 1 0 67804 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_738
timestamp 1704896540
transform 1 0 68908 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141_750
timestamp 1704896540
transform 1 0 70012 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_754
timestamp 1704896540
transform 1 0 70380 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_756
timestamp 1704896540
transform 1 0 70564 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_768
timestamp 1704896540
transform 1 0 71668 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_780
timestamp 1704896540
transform 1 0 72772 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141_792
timestamp 1704896540
transform 1 0 73876 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_800
timestamp 1704896540
transform 1 0 74612 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_702
timestamp 1704896540
transform 1 0 65596 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_714
timestamp 1704896540
transform 1 0 66700 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_726
timestamp 1704896540
transform 1 0 67804 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_728
timestamp 1704896540
transform 1 0 67988 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_740
timestamp 1704896540
transform 1 0 69092 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_752
timestamp 1704896540
transform 1 0 70196 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_764
timestamp 1704896540
transform 1 0 71300 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_142_776
timestamp 1704896540
transform 1 0 72404 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_782
timestamp 1704896540
transform 1 0 72956 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_784
timestamp 1704896540
transform 1 0 73140 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142_796
timestamp 1704896540
transform 1 0 74244 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_800
timestamp 1704896540
transform 1 0 74612 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_702
timestamp 1704896540
transform 1 0 65596 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_714
timestamp 1704896540
transform 1 0 66700 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_726
timestamp 1704896540
transform 1 0 67804 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_738
timestamp 1704896540
transform 1 0 68908 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143_750
timestamp 1704896540
transform 1 0 70012 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_754
timestamp 1704896540
transform 1 0 70380 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_756
timestamp 1704896540
transform 1 0 70564 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_768
timestamp 1704896540
transform 1 0 71668 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_780
timestamp 1704896540
transform 1 0 72772 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_143_792
timestamp 1704896540
transform 1 0 73876 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_800
timestamp 1704896540
transform 1 0 74612 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_702
timestamp 1704896540
transform 1 0 65596 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_714
timestamp 1704896540
transform 1 0 66700 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_726
timestamp 1704896540
transform 1 0 67804 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_728
timestamp 1704896540
transform 1 0 67988 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_740
timestamp 1704896540
transform 1 0 69092 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_752
timestamp 1704896540
transform 1 0 70196 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_764
timestamp 1704896540
transform 1 0 71300 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144_776
timestamp 1704896540
transform 1 0 72404 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_782
timestamp 1704896540
transform 1 0 72956 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_784
timestamp 1704896540
transform 1 0 73140 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144_796
timestamp 1704896540
transform 1 0 74244 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_800
timestamp 1704896540
transform 1 0 74612 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_702
timestamp 1704896540
transform 1 0 65596 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_714
timestamp 1704896540
transform 1 0 66700 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_726
timestamp 1704896540
transform 1 0 67804 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_738
timestamp 1704896540
transform 1 0 68908 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145_750
timestamp 1704896540
transform 1 0 70012 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_754
timestamp 1704896540
transform 1 0 70380 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_756
timestamp 1704896540
transform 1 0 70564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_768
timestamp 1704896540
transform 1 0 71668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_780
timestamp 1704896540
transform 1 0 72772 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145_792
timestamp 1704896540
transform 1 0 73876 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_800
timestamp 1704896540
transform 1 0 74612 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_702
timestamp 1704896540
transform 1 0 65596 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_714
timestamp 1704896540
transform 1 0 66700 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_726
timestamp 1704896540
transform 1 0 67804 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_728
timestamp 1704896540
transform 1 0 67988 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_740
timestamp 1704896540
transform 1 0 69092 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_752
timestamp 1704896540
transform 1 0 70196 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_764
timestamp 1704896540
transform 1 0 71300 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146_776
timestamp 1704896540
transform 1 0 72404 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_782
timestamp 1704896540
transform 1 0 72956 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_784
timestamp 1704896540
transform 1 0 73140 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146_796
timestamp 1704896540
transform 1 0 74244 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_800
timestamp 1704896540
transform 1 0 74612 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_702
timestamp 1704896540
transform 1 0 65596 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_714
timestamp 1704896540
transform 1 0 66700 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_726
timestamp 1704896540
transform 1 0 67804 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_738
timestamp 1704896540
transform 1 0 68908 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147_750
timestamp 1704896540
transform 1 0 70012 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_754
timestamp 1704896540
transform 1 0 70380 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_756
timestamp 1704896540
transform 1 0 70564 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_768
timestamp 1704896540
transform 1 0 71668 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_780
timestamp 1704896540
transform 1 0 72772 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147_792
timestamp 1704896540
transform 1 0 73876 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_800
timestamp 1704896540
transform 1 0 74612 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_702
timestamp 1704896540
transform 1 0 65596 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_714
timestamp 1704896540
transform 1 0 66700 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_726
timestamp 1704896540
transform 1 0 67804 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_728
timestamp 1704896540
transform 1 0 67988 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_740
timestamp 1704896540
transform 1 0 69092 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_752
timestamp 1704896540
transform 1 0 70196 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_764
timestamp 1704896540
transform 1 0 71300 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_148_776
timestamp 1704896540
transform 1 0 72404 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_782
timestamp 1704896540
transform 1 0 72956 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_784
timestamp 1704896540
transform 1 0 73140 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148_796
timestamp 1704896540
transform 1 0 74244 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_800
timestamp 1704896540
transform 1 0 74612 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_702
timestamp 1704896540
transform 1 0 65596 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_714
timestamp 1704896540
transform 1 0 66700 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_726
timestamp 1704896540
transform 1 0 67804 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_738
timestamp 1704896540
transform 1 0 68908 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149_750
timestamp 1704896540
transform 1 0 70012 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_754
timestamp 1704896540
transform 1 0 70380 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_756
timestamp 1704896540
transform 1 0 70564 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_768
timestamp 1704896540
transform 1 0 71668 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_780
timestamp 1704896540
transform 1 0 72772 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_149_792
timestamp 1704896540
transform 1 0 73876 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_800
timestamp 1704896540
transform 1 0 74612 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_702
timestamp 1704896540
transform 1 0 65596 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_714
timestamp 1704896540
transform 1 0 66700 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_726
timestamp 1704896540
transform 1 0 67804 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_728
timestamp 1704896540
transform 1 0 67988 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_740
timestamp 1704896540
transform 1 0 69092 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_752
timestamp 1704896540
transform 1 0 70196 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_764
timestamp 1704896540
transform 1 0 71300 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_150_776
timestamp 1704896540
transform 1 0 72404 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_782
timestamp 1704896540
transform 1 0 72956 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_784
timestamp 1704896540
transform 1 0 73140 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150_796
timestamp 1704896540
transform 1 0 74244 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_800
timestamp 1704896540
transform 1 0 74612 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_702
timestamp 1704896540
transform 1 0 65596 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_714
timestamp 1704896540
transform 1 0 66700 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_726
timestamp 1704896540
transform 1 0 67804 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_738
timestamp 1704896540
transform 1 0 68908 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151_750
timestamp 1704896540
transform 1 0 70012 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_754
timestamp 1704896540
transform 1 0 70380 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_756
timestamp 1704896540
transform 1 0 70564 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_768
timestamp 1704896540
transform 1 0 71668 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_780
timestamp 1704896540
transform 1 0 72772 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151_792
timestamp 1704896540
transform 1 0 73876 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_800
timestamp 1704896540
transform 1 0 74612 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_702
timestamp 1704896540
transform 1 0 65596 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_714
timestamp 1704896540
transform 1 0 66700 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_726
timestamp 1704896540
transform 1 0 67804 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_728
timestamp 1704896540
transform 1 0 67988 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_740
timestamp 1704896540
transform 1 0 69092 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_752
timestamp 1704896540
transform 1 0 70196 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_764
timestamp 1704896540
transform 1 0 71300 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_152_776
timestamp 1704896540
transform 1 0 72404 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_782
timestamp 1704896540
transform 1 0 72956 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_784
timestamp 1704896540
transform 1 0 73140 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152_796
timestamp 1704896540
transform 1 0 74244 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_800
timestamp 1704896540
transform 1 0 74612 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_702
timestamp 1704896540
transform 1 0 65596 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_714
timestamp 1704896540
transform 1 0 66700 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_726
timestamp 1704896540
transform 1 0 67804 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_738
timestamp 1704896540
transform 1 0 68908 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153_750
timestamp 1704896540
transform 1 0 70012 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_754
timestamp 1704896540
transform 1 0 70380 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_756
timestamp 1704896540
transform 1 0 70564 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_768
timestamp 1704896540
transform 1 0 71668 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_780
timestamp 1704896540
transform 1 0 72772 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153_792
timestamp 1704896540
transform 1 0 73876 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_800
timestamp 1704896540
transform 1 0 74612 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_702
timestamp 1704896540
transform 1 0 65596 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_714
timestamp 1704896540
transform 1 0 66700 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_726
timestamp 1704896540
transform 1 0 67804 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_728
timestamp 1704896540
transform 1 0 67988 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_740
timestamp 1704896540
transform 1 0 69092 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_752
timestamp 1704896540
transform 1 0 70196 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_764
timestamp 1704896540
transform 1 0 71300 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154_776
timestamp 1704896540
transform 1 0 72404 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_782
timestamp 1704896540
transform 1 0 72956 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_784
timestamp 1704896540
transform 1 0 73140 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154_796
timestamp 1704896540
transform 1 0 74244 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_800
timestamp 1704896540
transform 1 0 74612 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_702
timestamp 1704896540
transform 1 0 65596 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_714
timestamp 1704896540
transform 1 0 66700 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_726
timestamp 1704896540
transform 1 0 67804 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_728
timestamp 1704896540
transform 1 0 67988 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_740
timestamp 1704896540
transform 1 0 69092 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_752
timestamp 1704896540
transform 1 0 70196 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_756
timestamp 1704896540
transform 1 0 70564 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_768
timestamp 1704896540
transform 1 0 71668 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_780
timestamp 1704896540
transform 1 0 72772 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_784
timestamp 1704896540
transform 1 0 73140 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_155_796
timestamp 1704896540
transform 1 0 74244 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_800
timestamp 1704896540
transform 1 0 74612 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 39836 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform 1 0 51244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 46092 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 55200 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 63756 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 66332 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 25208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform 1 0 44436 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform 1 0 21988 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform 1 0 43332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform 1 0 65964 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 66332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform 1 0 37444 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform 1 0 50416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 67988 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 66332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 45632 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform 1 0 54096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform 1 0 41952 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform 1 0 17480 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform 1 0 41216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 70012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform 1 0 36156 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform 1 0 49128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 44528 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform 1 0 53360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform 1 0 70932 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform 1 0 33948 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform 1 0 48944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 73968 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 68724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform 1 0 41032 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform 1 0 52624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform 1 0 32476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform 1 0 48208 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform 1 0 47472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform 1 0 28980 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform 1 0 47472 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform 1 0 53268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 66332 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform 1 0 51152 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 66332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform 1 0 49404 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 66332 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform -1 0 49680 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 66332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform 1 0 54372 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 66332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 57408 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 66332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform 1 0 59156 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 66332 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform 1 0 57776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform -1 0 66332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform -1 0 35972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 66332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 62560 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 66332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 27416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform 1 0 45356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform 1 0 62928 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 66332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform -1 0 66332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform 1 0 31188 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 66332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform 1 0 46368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform 1 0 26036 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform 1 0 45632 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform 1 0 44896 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 23184 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform 1 0 43792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform 1 0 19872 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform 1 0 17572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform 1 0 40388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold86 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 42964 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform 1 0 19136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold89
timestamp 1704896540
transform 1 0 42320 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold92
timestamp 1704896540
transform 1 0 65596 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold95
timestamp 1704896540
transform 1 0 65596 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform 1 0 24564 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform 1 0 43700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform -1 0 46184 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform -1 0 35880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform 1 0 29716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform 1 0 15732 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform -1 0 46920 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform -1 0 47104 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform -1 0 41952 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform -1 0 40572 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 37260 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform 1 0 34868 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform 1 0 33212 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1704896540
transform -1 0 33212 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1704896540
transform 1 0 29716 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1704896540
transform -1 0 54832 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1704896540
transform -1 0 52256 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1704896540
transform -1 0 30176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1704896540
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1704896540
transform 1 0 47380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1704896540
transform 1 0 54096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1704896540
transform -1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1704896540
transform -1 0 60076 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1704896540
transform 1 0 55476 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1704896540
transform -1 0 65136 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1704896540
transform 1 0 57316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1704896540
transform -1 0 28244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1704896540
transform 1 0 60444 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1704896540
transform -1 0 23920 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1704896540
transform 1 0 62284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1704896540
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1704896540
transform -1 0 68816 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1704896540
transform -1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1704896540
transform -1 0 19136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1704896540
transform 1 0 69552 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1704896540
transform 1 0 70656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1704896540
transform 1 0 72312 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1704896540
transform -1 0 36708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1704896540
transform 1 0 32292 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1704896540
transform -1 0 32476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1704896540
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1704896540
transform 1 0 27140 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1704896540
transform -1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1704896540
transform 1 0 23460 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1704896540
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1704896540
transform 1 0 16744 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform -1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1704896540
transform -1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 44528 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 47104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1704896540
transform -1 0 20240 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1704896540
transform -1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1704896540
transform -1 0 25300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1704896540
transform 1 0 26864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1704896540
transform -1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1704896540
transform -1 0 28980 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1704896540
transform 1 0 32016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1704896540
transform -1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1704896540
transform -1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform 1 0 16192 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input15
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1704896540
transform 1 0 38180 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1704896540
transform -1 0 39652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 41768 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1704896540
transform -1 0 42780 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1704896540
transform -1 0 44804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1704896540
transform 1 0 46920 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1704896540
transform -1 0 47380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1704896540
transform 1 0 50140 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1704896540
transform 1 0 51888 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1704896540
transform 1 0 54096 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1704896540
transform -1 0 19780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1704896540
transform 1 0 55200 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1704896540
transform -1 0 56304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1704896540
transform 1 0 58512 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1704896540
transform 1 0 59892 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1704896540
transform -1 0 61180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1704896540
transform -1 0 63572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1704896540
transform 1 0 65504 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1704896540
transform 1 0 66700 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1704896540
transform -1 0 67804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1704896540
transform -1 0 69460 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input37
timestamp 1704896540
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input38
timestamp 1704896540
transform 1 0 71668 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input39
timestamp 1704896540
transform -1 0 73140 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input40
timestamp 1704896540
transform -1 0 25852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1704896540
transform -1 0 27876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1704896540
transform -1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1704896540
transform -1 0 31740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1704896540
transform -1 0 33120 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1704896540
transform -1 0 34684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1704896540
transform -1 0 36432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input47
timestamp 1704896540
transform 1 0 19780 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input48
timestamp 1704896540
transform 1 0 21988 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input49
timestamp 1704896540
transform 1 0 24196 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input50
timestamp 1704896540
transform 1 0 26864 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1704896540
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18032 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1704896540
transform -1 0 5152 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1704896540
transform -1 0 18032 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1704896540
transform -1 0 21528 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1704896540
transform 1 0 37996 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1704896540
transform 1 0 39744 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1704896540
transform 1 0 42320 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1704896540
transform 1 0 42964 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1704896540
transform 1 0 44896 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1704896540
transform 1 0 47472 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1704896540
transform 1 0 47932 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1704896540
transform 1 0 50048 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1704896540
transform 1 0 52624 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1704896540
transform 1 0 52900 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1704896540
transform -1 0 22908 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1704896540
transform 1 0 55200 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1704896540
transform 1 0 56212 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1704896540
transform 1 0 57868 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1704896540
transform 1 0 60352 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1704896540
transform 1 0 61180 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1704896540
transform 1 0 62928 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1704896540
transform 1 0 64492 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1704896540
transform 1 0 66148 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1704896540
transform 1 0 68080 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1704896540
transform 1 0 69460 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1704896540
transform -1 0 24196 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1704896540
transform 1 0 71116 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1704896540
transform 1 0 73232 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1704896540
transform -1 0 26772 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1704896540
transform 1 0 27876 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1704896540
transform 1 0 29716 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1704896540
transform 1 0 30452 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1704896540
transform 1 0 33028 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1704896540
transform 1 0 34684 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1704896540
transform 1 0 35604 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_0
timestamp 1704896540
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_9
timestamp 1704896540
transform -1 0 74980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_1
timestamp 1704896540
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_10
timestamp 1704896540
transform -1 0 74980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_2
timestamp 1704896540
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_11
timestamp 1704896540
transform -1 0 74980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_3
timestamp 1704896540
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_12
timestamp 1704896540
transform -1 0 74980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_4
timestamp 1704896540
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_13
timestamp 1704896540
transform -1 0 74980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_5
timestamp 1704896540
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_14
timestamp 1704896540
transform -1 0 74980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_6
timestamp 1704896540
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_15
timestamp 1704896540
transform -1 0 74980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_7
timestamp 1704896540
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_16
timestamp 1704896540
transform -1 0 74980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_8
timestamp 1704896540
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_17
timestamp 1704896540
transform -1 0 74980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_311
timestamp 1704896540
transform 1 0 65320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_164
timestamp 1704896540
transform -1 0 74980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_165
timestamp 1704896540
transform 1 0 65320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_18
timestamp 1704896540
transform -1 0 74980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_166
timestamp 1704896540
transform 1 0 65320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_19
timestamp 1704896540
transform -1 0 74980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_167
timestamp 1704896540
transform 1 0 65320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_20
timestamp 1704896540
transform -1 0 74980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_168
timestamp 1704896540
transform 1 0 65320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_21
timestamp 1704896540
transform -1 0 74980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_169
timestamp 1704896540
transform 1 0 65320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_22
timestamp 1704896540
transform -1 0 74980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_170
timestamp 1704896540
transform 1 0 65320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_23
timestamp 1704896540
transform -1 0 74980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_171
timestamp 1704896540
transform 1 0 65320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_24
timestamp 1704896540
transform -1 0 74980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_172
timestamp 1704896540
transform 1 0 65320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_25
timestamp 1704896540
transform -1 0 74980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_173
timestamp 1704896540
transform 1 0 65320 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_26
timestamp 1704896540
transform -1 0 74980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_174
timestamp 1704896540
transform 1 0 65320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_27
timestamp 1704896540
transform -1 0 74980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_175
timestamp 1704896540
transform 1 0 65320 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_28
timestamp 1704896540
transform -1 0 74980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_176
timestamp 1704896540
transform 1 0 65320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_29
timestamp 1704896540
transform -1 0 74980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_177
timestamp 1704896540
transform 1 0 65320 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_30
timestamp 1704896540
transform -1 0 74980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_178
timestamp 1704896540
transform 1 0 65320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_31
timestamp 1704896540
transform -1 0 74980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_179
timestamp 1704896540
transform 1 0 65320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_32
timestamp 1704896540
transform -1 0 74980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_180
timestamp 1704896540
transform 1 0 65320 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_33
timestamp 1704896540
transform -1 0 74980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_181
timestamp 1704896540
transform 1 0 65320 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_34
timestamp 1704896540
transform -1 0 74980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_182
timestamp 1704896540
transform 1 0 65320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_35
timestamp 1704896540
transform -1 0 74980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_183
timestamp 1704896540
transform 1 0 65320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_36
timestamp 1704896540
transform -1 0 74980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_184
timestamp 1704896540
transform 1 0 65320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_37
timestamp 1704896540
transform -1 0 74980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_185
timestamp 1704896540
transform 1 0 65320 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_38
timestamp 1704896540
transform -1 0 74980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_186
timestamp 1704896540
transform 1 0 65320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_39
timestamp 1704896540
transform -1 0 74980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_187
timestamp 1704896540
transform 1 0 65320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_40
timestamp 1704896540
transform -1 0 74980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_188
timestamp 1704896540
transform 1 0 65320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_41
timestamp 1704896540
transform -1 0 74980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_189
timestamp 1704896540
transform 1 0 65320 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_42
timestamp 1704896540
transform -1 0 74980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_190
timestamp 1704896540
transform 1 0 65320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_43
timestamp 1704896540
transform -1 0 74980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_191
timestamp 1704896540
transform 1 0 65320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_44
timestamp 1704896540
transform -1 0 74980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_192
timestamp 1704896540
transform 1 0 65320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_45
timestamp 1704896540
transform -1 0 74980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_193
timestamp 1704896540
transform 1 0 65320 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_46
timestamp 1704896540
transform -1 0 74980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_194
timestamp 1704896540
transform 1 0 65320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_47
timestamp 1704896540
transform -1 0 74980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_195
timestamp 1704896540
transform 1 0 65320 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_48
timestamp 1704896540
transform -1 0 74980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_196
timestamp 1704896540
transform 1 0 65320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_49
timestamp 1704896540
transform -1 0 74980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_197
timestamp 1704896540
transform 1 0 65320 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_50
timestamp 1704896540
transform -1 0 74980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_198
timestamp 1704896540
transform 1 0 65320 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_51
timestamp 1704896540
transform -1 0 74980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_199
timestamp 1704896540
transform 1 0 65320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_52
timestamp 1704896540
transform -1 0 74980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_200
timestamp 1704896540
transform 1 0 65320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_53
timestamp 1704896540
transform -1 0 74980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_201
timestamp 1704896540
transform 1 0 65320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_54
timestamp 1704896540
transform -1 0 74980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_202
timestamp 1704896540
transform 1 0 65320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_55
timestamp 1704896540
transform -1 0 74980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_203
timestamp 1704896540
transform 1 0 65320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_56
timestamp 1704896540
transform -1 0 74980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_204
timestamp 1704896540
transform 1 0 65320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_57
timestamp 1704896540
transform -1 0 74980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_205
timestamp 1704896540
transform 1 0 65320 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_58
timestamp 1704896540
transform -1 0 74980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_206
timestamp 1704896540
transform 1 0 65320 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_59
timestamp 1704896540
transform -1 0 74980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_207
timestamp 1704896540
transform 1 0 65320 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_60
timestamp 1704896540
transform -1 0 74980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_208
timestamp 1704896540
transform 1 0 65320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_61
timestamp 1704896540
transform -1 0 74980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_209
timestamp 1704896540
transform 1 0 65320 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_62
timestamp 1704896540
transform -1 0 74980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_210
timestamp 1704896540
transform 1 0 65320 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_63
timestamp 1704896540
transform -1 0 74980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_211
timestamp 1704896540
transform 1 0 65320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_64
timestamp 1704896540
transform -1 0 74980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_212
timestamp 1704896540
transform 1 0 65320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_65
timestamp 1704896540
transform -1 0 74980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_213
timestamp 1704896540
transform 1 0 65320 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_66
timestamp 1704896540
transform -1 0 74980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_214
timestamp 1704896540
transform 1 0 65320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_67
timestamp 1704896540
transform -1 0 74980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_215
timestamp 1704896540
transform 1 0 65320 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_68
timestamp 1704896540
transform -1 0 74980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_216
timestamp 1704896540
transform 1 0 65320 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_69
timestamp 1704896540
transform -1 0 74980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_217
timestamp 1704896540
transform 1 0 65320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_70
timestamp 1704896540
transform -1 0 74980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_218
timestamp 1704896540
transform 1 0 65320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_71
timestamp 1704896540
transform -1 0 74980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_219
timestamp 1704896540
transform 1 0 65320 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_72
timestamp 1704896540
transform -1 0 74980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_220
timestamp 1704896540
transform 1 0 65320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_73
timestamp 1704896540
transform -1 0 74980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_221
timestamp 1704896540
transform 1 0 65320 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_74
timestamp 1704896540
transform -1 0 74980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_222
timestamp 1704896540
transform 1 0 65320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_75
timestamp 1704896540
transform -1 0 74980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_223
timestamp 1704896540
transform 1 0 65320 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_76
timestamp 1704896540
transform -1 0 74980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_224
timestamp 1704896540
transform 1 0 65320 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_77
timestamp 1704896540
transform -1 0 74980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_225
timestamp 1704896540
transform 1 0 65320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_78
timestamp 1704896540
transform -1 0 74980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_226
timestamp 1704896540
transform 1 0 65320 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_79
timestamp 1704896540
transform -1 0 74980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_227
timestamp 1704896540
transform 1 0 65320 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_80
timestamp 1704896540
transform -1 0 74980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_228
timestamp 1704896540
transform 1 0 65320 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_81
timestamp 1704896540
transform -1 0 74980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_229
timestamp 1704896540
transform 1 0 65320 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_82
timestamp 1704896540
transform -1 0 74980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_230
timestamp 1704896540
transform 1 0 65320 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_83
timestamp 1704896540
transform -1 0 74980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_231
timestamp 1704896540
transform 1 0 65320 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_84
timestamp 1704896540
transform -1 0 74980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_232
timestamp 1704896540
transform 1 0 65320 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_85
timestamp 1704896540
transform -1 0 74980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_233
timestamp 1704896540
transform 1 0 65320 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_86
timestamp 1704896540
transform -1 0 74980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_234
timestamp 1704896540
transform 1 0 65320 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_87
timestamp 1704896540
transform -1 0 74980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_235
timestamp 1704896540
transform 1 0 65320 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_88
timestamp 1704896540
transform -1 0 74980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_236
timestamp 1704896540
transform 1 0 65320 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_89
timestamp 1704896540
transform -1 0 74980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_237
timestamp 1704896540
transform 1 0 65320 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_90
timestamp 1704896540
transform -1 0 74980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_238
timestamp 1704896540
transform 1 0 65320 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_91
timestamp 1704896540
transform -1 0 74980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_239
timestamp 1704896540
transform 1 0 65320 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_92
timestamp 1704896540
transform -1 0 74980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_240
timestamp 1704896540
transform 1 0 65320 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_93
timestamp 1704896540
transform -1 0 74980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_241
timestamp 1704896540
transform 1 0 65320 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_94
timestamp 1704896540
transform -1 0 74980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_242
timestamp 1704896540
transform 1 0 65320 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_95
timestamp 1704896540
transform -1 0 74980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_243
timestamp 1704896540
transform 1 0 65320 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_96
timestamp 1704896540
transform -1 0 74980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_244
timestamp 1704896540
transform 1 0 65320 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_97
timestamp 1704896540
transform -1 0 74980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_245
timestamp 1704896540
transform 1 0 65320 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_98
timestamp 1704896540
transform -1 0 74980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_246
timestamp 1704896540
transform 1 0 65320 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_99
timestamp 1704896540
transform -1 0 74980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_247
timestamp 1704896540
transform 1 0 65320 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_100
timestamp 1704896540
transform -1 0 74980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_248
timestamp 1704896540
transform 1 0 65320 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_101
timestamp 1704896540
transform -1 0 74980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_249
timestamp 1704896540
transform 1 0 65320 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_102
timestamp 1704896540
transform -1 0 74980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_250
timestamp 1704896540
transform 1 0 65320 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_103
timestamp 1704896540
transform -1 0 74980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_251
timestamp 1704896540
transform 1 0 65320 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_104
timestamp 1704896540
transform -1 0 74980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_252
timestamp 1704896540
transform 1 0 65320 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_105
timestamp 1704896540
transform -1 0 74980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_253
timestamp 1704896540
transform 1 0 65320 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_106
timestamp 1704896540
transform -1 0 74980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_254
timestamp 1704896540
transform 1 0 65320 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_107
timestamp 1704896540
transform -1 0 74980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_255
timestamp 1704896540
transform 1 0 65320 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_108
timestamp 1704896540
transform -1 0 74980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_256
timestamp 1704896540
transform 1 0 65320 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_109
timestamp 1704896540
transform -1 0 74980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_257
timestamp 1704896540
transform 1 0 65320 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_110
timestamp 1704896540
transform -1 0 74980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_258
timestamp 1704896540
transform 1 0 65320 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_111
timestamp 1704896540
transform -1 0 74980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_259
timestamp 1704896540
transform 1 0 65320 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_112
timestamp 1704896540
transform -1 0 74980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_260
timestamp 1704896540
transform 1 0 65320 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_113
timestamp 1704896540
transform -1 0 74980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_261
timestamp 1704896540
transform 1 0 65320 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_114
timestamp 1704896540
transform -1 0 74980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_262
timestamp 1704896540
transform 1 0 65320 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_115
timestamp 1704896540
transform -1 0 74980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_263
timestamp 1704896540
transform 1 0 65320 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_116
timestamp 1704896540
transform -1 0 74980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_264
timestamp 1704896540
transform 1 0 65320 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_117
timestamp 1704896540
transform -1 0 74980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_265
timestamp 1704896540
transform 1 0 65320 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_118
timestamp 1704896540
transform -1 0 74980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_266
timestamp 1704896540
transform 1 0 65320 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_119
timestamp 1704896540
transform -1 0 74980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_267
timestamp 1704896540
transform 1 0 65320 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_120
timestamp 1704896540
transform -1 0 74980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_268
timestamp 1704896540
transform 1 0 65320 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_121
timestamp 1704896540
transform -1 0 74980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_269
timestamp 1704896540
transform 1 0 65320 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_122
timestamp 1704896540
transform -1 0 74980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_270
timestamp 1704896540
transform 1 0 65320 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_123
timestamp 1704896540
transform -1 0 74980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_271
timestamp 1704896540
transform 1 0 65320 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_124
timestamp 1704896540
transform -1 0 74980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Left_272
timestamp 1704896540
transform 1 0 65320 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Right_125
timestamp 1704896540
transform -1 0 74980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Left_273
timestamp 1704896540
transform 1 0 65320 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Right_126
timestamp 1704896540
transform -1 0 74980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Left_274
timestamp 1704896540
transform 1 0 65320 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Right_127
timestamp 1704896540
transform -1 0 74980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Left_275
timestamp 1704896540
transform 1 0 65320 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Right_128
timestamp 1704896540
transform -1 0 74980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_276
timestamp 1704896540
transform 1 0 65320 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_129
timestamp 1704896540
transform -1 0 74980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_277
timestamp 1704896540
transform 1 0 65320 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_130
timestamp 1704896540
transform -1 0 74980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_278
timestamp 1704896540
transform 1 0 65320 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_131
timestamp 1704896540
transform -1 0 74980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_279
timestamp 1704896540
transform 1 0 65320 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_132
timestamp 1704896540
transform -1 0 74980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_280
timestamp 1704896540
transform 1 0 65320 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_133
timestamp 1704896540
transform -1 0 74980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_281
timestamp 1704896540
transform 1 0 65320 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_134
timestamp 1704896540
transform -1 0 74980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_282
timestamp 1704896540
transform 1 0 65320 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_135
timestamp 1704896540
transform -1 0 74980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_283
timestamp 1704896540
transform 1 0 65320 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_136
timestamp 1704896540
transform -1 0 74980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_284
timestamp 1704896540
transform 1 0 65320 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_137
timestamp 1704896540
transform -1 0 74980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_285
timestamp 1704896540
transform 1 0 65320 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_138
timestamp 1704896540
transform -1 0 74980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_286
timestamp 1704896540
transform 1 0 65320 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_139
timestamp 1704896540
transform -1 0 74980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_287
timestamp 1704896540
transform 1 0 65320 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_140
timestamp 1704896540
transform -1 0 74980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_288
timestamp 1704896540
transform 1 0 65320 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_141
timestamp 1704896540
transform -1 0 74980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_289
timestamp 1704896540
transform 1 0 65320 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_142
timestamp 1704896540
transform -1 0 74980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_290
timestamp 1704896540
transform 1 0 65320 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_143
timestamp 1704896540
transform -1 0 74980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_291
timestamp 1704896540
transform 1 0 65320 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_144
timestamp 1704896540
transform -1 0 74980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_292
timestamp 1704896540
transform 1 0 65320 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_145
timestamp 1704896540
transform -1 0 74980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_293
timestamp 1704896540
transform 1 0 65320 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_146
timestamp 1704896540
transform -1 0 74980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_294
timestamp 1704896540
transform 1 0 65320 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_147
timestamp 1704896540
transform -1 0 74980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_295
timestamp 1704896540
transform 1 0 65320 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_148
timestamp 1704896540
transform -1 0 74980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_296
timestamp 1704896540
transform 1 0 65320 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_149
timestamp 1704896540
transform -1 0 74980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_297
timestamp 1704896540
transform 1 0 65320 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_150
timestamp 1704896540
transform -1 0 74980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_298
timestamp 1704896540
transform 1 0 65320 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_151
timestamp 1704896540
transform -1 0 74980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_299
timestamp 1704896540
transform 1 0 65320 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_152
timestamp 1704896540
transform -1 0 74980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_300
timestamp 1704896540
transform 1 0 65320 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_153
timestamp 1704896540
transform -1 0 74980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_301
timestamp 1704896540
transform 1 0 65320 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_154
timestamp 1704896540
transform -1 0 74980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_302
timestamp 1704896540
transform 1 0 65320 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_155
timestamp 1704896540
transform -1 0 74980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_303
timestamp 1704896540
transform 1 0 65320 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_156
timestamp 1704896540
transform -1 0 74980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_304
timestamp 1704896540
transform 1 0 65320 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_157
timestamp 1704896540
transform -1 0 74980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_305
timestamp 1704896540
transform 1 0 65320 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_158
timestamp 1704896540
transform -1 0 74980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_306
timestamp 1704896540
transform 1 0 65320 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_159
timestamp 1704896540
transform -1 0 74980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_307
timestamp 1704896540
transform 1 0 65320 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_160
timestamp 1704896540
transform -1 0 74980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_308
timestamp 1704896540
transform 1 0 65320 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_161
timestamp 1704896540
transform -1 0 74980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_309
timestamp 1704896540
transform 1 0 65320 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_162
timestamp 1704896540
transform -1 0 74980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_310
timestamp 1704896540
transform 1 0 65320 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_163
timestamp 1704896540
transform -1 0 74980 0 -1 85952
box -38 -48 314 592
use EFSRAM_1024x32_wrapper  SRAM_0
timestamp 0
transform 0 -1 63283 1 0 8000
box 0 -40 77574 61263
use sky130_fd_sc_hd__conb_1  SRAM_0_87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 65872 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_88
timestamp 1704896540
transform -1 0 65872 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_89
timestamp 1704896540
transform -1 0 65872 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_90
timestamp 1704896540
transform -1 0 65872 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_91
timestamp 1704896540
transform -1 0 65872 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_92
timestamp 1704896540
transform -1 0 66148 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_93
timestamp 1704896540
transform -1 0 65872 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_94
timestamp 1704896540
transform 1 0 65596 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_95
timestamp 1704896540
transform 1 0 65872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_312 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_313
timestamp 1704896540
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_314
timestamp 1704896540
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_315
timestamp 1704896540
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_316
timestamp 1704896540
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_317
timestamp 1704896540
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_318
timestamp 1704896540
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_319
timestamp 1704896540
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_320
timestamp 1704896540
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_321
timestamp 1704896540
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_322
timestamp 1704896540
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_323
timestamp 1704896540
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_324
timestamp 1704896540
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_325
timestamp 1704896540
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_326
timestamp 1704896540
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_327
timestamp 1704896540
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_328
timestamp 1704896540
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_329
timestamp 1704896540
transform 1 0 47380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_330
timestamp 1704896540
transform 1 0 49956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_331
timestamp 1704896540
transform 1 0 52532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_332
timestamp 1704896540
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_333
timestamp 1704896540
transform 1 0 57684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_334
timestamp 1704896540
transform 1 0 60260 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_335
timestamp 1704896540
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_336
timestamp 1704896540
transform 1 0 65412 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_337
timestamp 1704896540
transform 1 0 67988 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_338
timestamp 1704896540
transform 1 0 70564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_339
timestamp 1704896540
transform 1 0 73140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_340
timestamp 1704896540
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_341
timestamp 1704896540
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_342
timestamp 1704896540
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_343
timestamp 1704896540
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_344
timestamp 1704896540
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_345
timestamp 1704896540
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_346
timestamp 1704896540
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_347
timestamp 1704896540
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_348
timestamp 1704896540
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_349
timestamp 1704896540
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_350
timestamp 1704896540
transform 1 0 57684 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_351
timestamp 1704896540
transform 1 0 62836 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_352
timestamp 1704896540
transform 1 0 67988 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_353
timestamp 1704896540
transform 1 0 73140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_354
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_355
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_356
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_357
timestamp 1704896540
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_358
timestamp 1704896540
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_359
timestamp 1704896540
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_360
timestamp 1704896540
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_361
timestamp 1704896540
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_362
timestamp 1704896540
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_363
timestamp 1704896540
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_364
timestamp 1704896540
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_365
timestamp 1704896540
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_366
timestamp 1704896540
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_367
timestamp 1704896540
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_368
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_369
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_370
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_371
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_372
timestamp 1704896540
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_373
timestamp 1704896540
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_374
timestamp 1704896540
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_375
timestamp 1704896540
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_376
timestamp 1704896540
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_377
timestamp 1704896540
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_378
timestamp 1704896540
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_379
timestamp 1704896540
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_380
timestamp 1704896540
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_381
timestamp 1704896540
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_382
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_383
timestamp 1704896540
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_384
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_385
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_386
timestamp 1704896540
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_387
timestamp 1704896540
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_388
timestamp 1704896540
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_389
timestamp 1704896540
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_390
timestamp 1704896540
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_391
timestamp 1704896540
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_392
timestamp 1704896540
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_393
timestamp 1704896540
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_394
timestamp 1704896540
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_395
timestamp 1704896540
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_396
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_397
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_398
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_399
timestamp 1704896540
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_400
timestamp 1704896540
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_401
timestamp 1704896540
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_402
timestamp 1704896540
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_403
timestamp 1704896540
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_404
timestamp 1704896540
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_405
timestamp 1704896540
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_406
timestamp 1704896540
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_407
timestamp 1704896540
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_408
timestamp 1704896540
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_409
timestamp 1704896540
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_410
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_411
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_412
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_413
timestamp 1704896540
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_414
timestamp 1704896540
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_415
timestamp 1704896540
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_416
timestamp 1704896540
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_417
timestamp 1704896540
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_418
timestamp 1704896540
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_419
timestamp 1704896540
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_420
timestamp 1704896540
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_421
timestamp 1704896540
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_422
timestamp 1704896540
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_423
timestamp 1704896540
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_424
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_425
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_426
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_427
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_428
timestamp 1704896540
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_429
timestamp 1704896540
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_430
timestamp 1704896540
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_431
timestamp 1704896540
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_432
timestamp 1704896540
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_433
timestamp 1704896540
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_434
timestamp 1704896540
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_435
timestamp 1704896540
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_436
timestamp 1704896540
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_437
timestamp 1704896540
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_438
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_439
timestamp 1704896540
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_440
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_441
timestamp 1704896540
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_442
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_443
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_444
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_445
timestamp 1704896540
transform 1 0 21620 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_446
timestamp 1704896540
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_447
timestamp 1704896540
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_448
timestamp 1704896540
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_449
timestamp 1704896540
transform 1 0 31924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_450
timestamp 1704896540
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_451
timestamp 1704896540
transform 1 0 37076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_452
timestamp 1704896540
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_453
timestamp 1704896540
transform 1 0 42228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_454
timestamp 1704896540
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_455
timestamp 1704896540
transform 1 0 47380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_456
timestamp 1704896540
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_457
timestamp 1704896540
transform 1 0 52532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_458
timestamp 1704896540
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_459
timestamp 1704896540
transform 1 0 57684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_460
timestamp 1704896540
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_461
timestamp 1704896540
transform 1 0 62836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_462
timestamp 1704896540
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_463
timestamp 1704896540
transform 1 0 67988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_464
timestamp 1704896540
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_465
timestamp 1704896540
transform 1 0 73140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_687
timestamp 1704896540
transform 1 0 70472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_466
timestamp 1704896540
transform 1 0 67896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_467
timestamp 1704896540
transform 1 0 73048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_468
timestamp 1704896540
transform 1 0 70472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_469
timestamp 1704896540
transform 1 0 67896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_470
timestamp 1704896540
transform 1 0 73048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_471
timestamp 1704896540
transform 1 0 70472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_472
timestamp 1704896540
transform 1 0 67896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_473
timestamp 1704896540
transform 1 0 73048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_474
timestamp 1704896540
transform 1 0 70472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_475
timestamp 1704896540
transform 1 0 67896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_476
timestamp 1704896540
transform 1 0 73048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_477
timestamp 1704896540
transform 1 0 70472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_478
timestamp 1704896540
transform 1 0 67896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_479
timestamp 1704896540
transform 1 0 73048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_480
timestamp 1704896540
transform 1 0 70472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_481
timestamp 1704896540
transform 1 0 67896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_482
timestamp 1704896540
transform 1 0 73048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_483
timestamp 1704896540
transform 1 0 70472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_484
timestamp 1704896540
transform 1 0 67896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_485
timestamp 1704896540
transform 1 0 73048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_486
timestamp 1704896540
transform 1 0 70472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_487
timestamp 1704896540
transform 1 0 67896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_488
timestamp 1704896540
transform 1 0 73048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_489
timestamp 1704896540
transform 1 0 70472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_490
timestamp 1704896540
transform 1 0 67896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_491
timestamp 1704896540
transform 1 0 73048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_492
timestamp 1704896540
transform 1 0 70472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_493
timestamp 1704896540
transform 1 0 67896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_494
timestamp 1704896540
transform 1 0 73048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_495
timestamp 1704896540
transform 1 0 70472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_496
timestamp 1704896540
transform 1 0 67896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_497
timestamp 1704896540
transform 1 0 73048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_498
timestamp 1704896540
transform 1 0 70472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_499
timestamp 1704896540
transform 1 0 67896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_500
timestamp 1704896540
transform 1 0 73048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_501
timestamp 1704896540
transform 1 0 70472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_502
timestamp 1704896540
transform 1 0 67896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_503
timestamp 1704896540
transform 1 0 73048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_504
timestamp 1704896540
transform 1 0 70472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_505
timestamp 1704896540
transform 1 0 67896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_506
timestamp 1704896540
transform 1 0 73048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_507
timestamp 1704896540
transform 1 0 70472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_508
timestamp 1704896540
transform 1 0 67896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_509
timestamp 1704896540
transform 1 0 73048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_510
timestamp 1704896540
transform 1 0 70472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_511
timestamp 1704896540
transform 1 0 67896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_512
timestamp 1704896540
transform 1 0 73048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_513
timestamp 1704896540
transform 1 0 70472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_514
timestamp 1704896540
transform 1 0 67896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_515
timestamp 1704896540
transform 1 0 73048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_516
timestamp 1704896540
transform 1 0 70472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_517
timestamp 1704896540
transform 1 0 67896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_518
timestamp 1704896540
transform 1 0 73048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_519
timestamp 1704896540
transform 1 0 70472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_520
timestamp 1704896540
transform 1 0 67896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_521
timestamp 1704896540
transform 1 0 73048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_522
timestamp 1704896540
transform 1 0 70472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_523
timestamp 1704896540
transform 1 0 67896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_524
timestamp 1704896540
transform 1 0 73048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_525
timestamp 1704896540
transform 1 0 70472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_526
timestamp 1704896540
transform 1 0 67896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_527
timestamp 1704896540
transform 1 0 73048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_528
timestamp 1704896540
transform 1 0 70472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_529
timestamp 1704896540
transform 1 0 67896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_530
timestamp 1704896540
transform 1 0 73048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_531
timestamp 1704896540
transform 1 0 70472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_532
timestamp 1704896540
transform 1 0 67896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_533
timestamp 1704896540
transform 1 0 73048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_534
timestamp 1704896540
transform 1 0 70472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_535
timestamp 1704896540
transform 1 0 67896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_536
timestamp 1704896540
transform 1 0 73048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_537
timestamp 1704896540
transform 1 0 70472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_538
timestamp 1704896540
transform 1 0 67896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_539
timestamp 1704896540
transform 1 0 73048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_540
timestamp 1704896540
transform 1 0 70472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_541
timestamp 1704896540
transform 1 0 67896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_542
timestamp 1704896540
transform 1 0 73048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_543
timestamp 1704896540
transform 1 0 70472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_544
timestamp 1704896540
transform 1 0 67896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_545
timestamp 1704896540
transform 1 0 73048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_546
timestamp 1704896540
transform 1 0 70472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_547
timestamp 1704896540
transform 1 0 67896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_548
timestamp 1704896540
transform 1 0 73048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_549
timestamp 1704896540
transform 1 0 70472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_550
timestamp 1704896540
transform 1 0 67896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_551
timestamp 1704896540
transform 1 0 73048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_552
timestamp 1704896540
transform 1 0 70472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_553
timestamp 1704896540
transform 1 0 67896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_554
timestamp 1704896540
transform 1 0 73048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_555
timestamp 1704896540
transform 1 0 70472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_556
timestamp 1704896540
transform 1 0 67896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_557
timestamp 1704896540
transform 1 0 73048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_558
timestamp 1704896540
transform 1 0 70472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_559
timestamp 1704896540
transform 1 0 67896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_560
timestamp 1704896540
transform 1 0 73048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_561
timestamp 1704896540
transform 1 0 70472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_562
timestamp 1704896540
transform 1 0 67896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_563
timestamp 1704896540
transform 1 0 73048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_564
timestamp 1704896540
transform 1 0 70472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_565
timestamp 1704896540
transform 1 0 67896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_566
timestamp 1704896540
transform 1 0 73048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_567
timestamp 1704896540
transform 1 0 70472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_568
timestamp 1704896540
transform 1 0 67896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_569
timestamp 1704896540
transform 1 0 73048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_570
timestamp 1704896540
transform 1 0 70472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_571
timestamp 1704896540
transform 1 0 67896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_572
timestamp 1704896540
transform 1 0 73048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_573
timestamp 1704896540
transform 1 0 70472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_574
timestamp 1704896540
transform 1 0 67896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_575
timestamp 1704896540
transform 1 0 73048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_576
timestamp 1704896540
transform 1 0 70472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_577
timestamp 1704896540
transform 1 0 67896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_578
timestamp 1704896540
transform 1 0 73048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_579
timestamp 1704896540
transform 1 0 70472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_580
timestamp 1704896540
transform 1 0 67896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_581
timestamp 1704896540
transform 1 0 73048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_582
timestamp 1704896540
transform 1 0 70472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_583
timestamp 1704896540
transform 1 0 67896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_584
timestamp 1704896540
transform 1 0 73048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_585
timestamp 1704896540
transform 1 0 70472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_586
timestamp 1704896540
transform 1 0 67896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_587
timestamp 1704896540
transform 1 0 73048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_588
timestamp 1704896540
transform 1 0 70472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_589
timestamp 1704896540
transform 1 0 67896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_590
timestamp 1704896540
transform 1 0 73048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_591
timestamp 1704896540
transform 1 0 70472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_592
timestamp 1704896540
transform 1 0 67896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_593
timestamp 1704896540
transform 1 0 73048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_594
timestamp 1704896540
transform 1 0 70472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_595
timestamp 1704896540
transform 1 0 67896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_596
timestamp 1704896540
transform 1 0 73048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_597
timestamp 1704896540
transform 1 0 70472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_598
timestamp 1704896540
transform 1 0 67896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_599
timestamp 1704896540
transform 1 0 73048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_600
timestamp 1704896540
transform 1 0 70472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_601
timestamp 1704896540
transform 1 0 67896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_602
timestamp 1704896540
transform 1 0 73048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_603
timestamp 1704896540
transform 1 0 70472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_604
timestamp 1704896540
transform 1 0 67896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_605
timestamp 1704896540
transform 1 0 73048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_606
timestamp 1704896540
transform 1 0 70472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_607
timestamp 1704896540
transform 1 0 67896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_608
timestamp 1704896540
transform 1 0 73048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_609
timestamp 1704896540
transform 1 0 70472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_610
timestamp 1704896540
transform 1 0 67896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_611
timestamp 1704896540
transform 1 0 73048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_612
timestamp 1704896540
transform 1 0 70472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_613
timestamp 1704896540
transform 1 0 67896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_614
timestamp 1704896540
transform 1 0 73048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_615
timestamp 1704896540
transform 1 0 70472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_616
timestamp 1704896540
transform 1 0 67896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_617
timestamp 1704896540
transform 1 0 73048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_618
timestamp 1704896540
transform 1 0 70472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_619
timestamp 1704896540
transform 1 0 67896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_620
timestamp 1704896540
transform 1 0 73048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_621
timestamp 1704896540
transform 1 0 70472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_622
timestamp 1704896540
transform 1 0 67896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_623
timestamp 1704896540
transform 1 0 73048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_624
timestamp 1704896540
transform 1 0 70472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_625
timestamp 1704896540
transform 1 0 67896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_626
timestamp 1704896540
transform 1 0 73048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_627
timestamp 1704896540
transform 1 0 70472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_628
timestamp 1704896540
transform 1 0 67896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_629
timestamp 1704896540
transform 1 0 73048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_630
timestamp 1704896540
transform 1 0 70472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_631
timestamp 1704896540
transform 1 0 67896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_632
timestamp 1704896540
transform 1 0 73048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_633
timestamp 1704896540
transform 1 0 70472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_634
timestamp 1704896540
transform 1 0 67896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_635
timestamp 1704896540
transform 1 0 73048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_636
timestamp 1704896540
transform 1 0 70472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_637
timestamp 1704896540
transform 1 0 67896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_638
timestamp 1704896540
transform 1 0 73048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_639
timestamp 1704896540
transform 1 0 70472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_640
timestamp 1704896540
transform 1 0 67896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_641
timestamp 1704896540
transform 1 0 73048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_642
timestamp 1704896540
transform 1 0 70472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_643
timestamp 1704896540
transform 1 0 67896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_644
timestamp 1704896540
transform 1 0 73048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_645
timestamp 1704896540
transform 1 0 70472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_646
timestamp 1704896540
transform 1 0 67896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_647
timestamp 1704896540
transform 1 0 73048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_648
timestamp 1704896540
transform 1 0 70472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_649
timestamp 1704896540
transform 1 0 67896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_650
timestamp 1704896540
transform 1 0 73048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_651
timestamp 1704896540
transform 1 0 70472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_652
timestamp 1704896540
transform 1 0 67896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_653
timestamp 1704896540
transform 1 0 73048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_654
timestamp 1704896540
transform 1 0 70472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_655
timestamp 1704896540
transform 1 0 67896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_656
timestamp 1704896540
transform 1 0 73048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_657
timestamp 1704896540
transform 1 0 70472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_658
timestamp 1704896540
transform 1 0 67896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_659
timestamp 1704896540
transform 1 0 73048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_660
timestamp 1704896540
transform 1 0 70472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_661
timestamp 1704896540
transform 1 0 67896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_662
timestamp 1704896540
transform 1 0 73048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_663
timestamp 1704896540
transform 1 0 70472 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_664
timestamp 1704896540
transform 1 0 67896 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_665
timestamp 1704896540
transform 1 0 73048 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_666
timestamp 1704896540
transform 1 0 70472 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_667
timestamp 1704896540
transform 1 0 67896 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_668
timestamp 1704896540
transform 1 0 73048 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_669
timestamp 1704896540
transform 1 0 70472 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_670
timestamp 1704896540
transform 1 0 67896 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_671
timestamp 1704896540
transform 1 0 73048 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_672
timestamp 1704896540
transform 1 0 70472 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_673
timestamp 1704896540
transform 1 0 67896 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_674
timestamp 1704896540
transform 1 0 73048 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_675
timestamp 1704896540
transform 1 0 70472 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_676
timestamp 1704896540
transform 1 0 67896 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_677
timestamp 1704896540
transform 1 0 73048 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_678
timestamp 1704896540
transform 1 0 70472 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_679
timestamp 1704896540
transform 1 0 67896 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_680
timestamp 1704896540
transform 1 0 73048 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_681
timestamp 1704896540
transform 1 0 70472 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_682
timestamp 1704896540
transform 1 0 67896 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_683
timestamp 1704896540
transform 1 0 73048 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_684
timestamp 1704896540
transform 1 0 67896 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_685
timestamp 1704896540
transform 1 0 70472 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_686
timestamp 1704896540
transform 1 0 73048 0 -1 85952
box -38 -48 130 592
<< labels >>
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 sram_selected
port 0 nsew signal tristate
flabel metal2 s 1836 1040 2188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 11836 1040 12188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 21836 1040 22188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 31836 1040 32188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 41836 1040 42188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 51836 1040 52188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 61836 1040 62188 7944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 71836 1040 72188 86000 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 1912 75028 2264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 11912 75028 12264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 21912 75028 22264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 31912 75028 32264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 41912 75028 42264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 51912 75028 52264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 61912 75028 62264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 71912 75028 72264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 81912 75028 82264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 86940 2322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 86940 8322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 86940 14322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 86940 20322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 86940 26322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 86940 32322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 86940 38322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 86940 44322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 86940 50322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 86940 56322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 86940 62322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 86940 68322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 86940 74322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 4188 1040 4540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 14188 1040 14540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 24188 1040 24540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 34188 1040 34540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 44188 1040 44540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 54188 1040 54540 7944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 64188 1040 64540 86000 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 74188 1040 74540 86000 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 4264 75028 4616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 14264 75028 14616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 24264 75028 24616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 34264 75028 34616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 44264 75028 44616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 54264 75028 54616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 64264 75028 64616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 74264 75028 74616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 84264 75028 84616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 0 5322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 0 5322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 86940 5322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 0 11322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 0 11322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 86940 11322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 0 17322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 0 17322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 86940 17322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 0 23322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 0 23322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 86940 23322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 0 29322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 0 29322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 86940 29322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 0 35322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 0 35322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 86940 35322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 0 41322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 0 41322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 86940 41322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 0 47322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 0 47322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 86940 47322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 0 53322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 0 53322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 86940 53322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 0 59322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 0 59322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 86940 59322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 0 65322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 0 65322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 86940 65322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 0 71322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 0 71322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 86940 71322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wb_clk_i
port 3 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wb_rst_i
port 4 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 5 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 6 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 7 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 8 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 9 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 10 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 11 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 12 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 13 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 14 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 15 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 16 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 17 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 18 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 19 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 20 nsew signal input
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 21 nsew signal input
flabel metal2 s 60002 0 60058 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 22 nsew signal input
flabel metal2 s 61658 0 61714 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 23 nsew signal input
flabel metal2 s 63314 0 63370 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 24 nsew signal input
flabel metal2 s 64970 0 65026 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 25 nsew signal input
flabel metal2 s 66626 0 66682 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 26 nsew signal input
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 27 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 28 nsew signal input
flabel metal2 s 69938 0 69994 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 29 nsew signal input
flabel metal2 s 71594 0 71650 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 30 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 31 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 32 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 33 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 34 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 35 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 36 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 37 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 38 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 39 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 40 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 41 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 42 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 43 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 44 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 45 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 46 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 47 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 48 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 49 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 50 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 51 nsew signal input
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 52 nsew signal input
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 53 nsew signal input
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 54 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 55 nsew signal input
flabel metal2 s 62210 0 62266 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 56 nsew signal input
flabel metal2 s 63866 0 63922 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 57 nsew signal input
flabel metal2 s 65522 0 65578 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 58 nsew signal input
flabel metal2 s 67178 0 67234 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 59 nsew signal input
flabel metal2 s 68834 0 68890 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 60 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 61 nsew signal input
flabel metal2 s 70490 0 70546 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 62 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 63 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 64 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 65 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 66 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 67 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 68 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 69 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 70 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 71 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 72 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 73 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 74 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 75 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 76 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 77 nsew signal tristate
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 78 nsew signal tristate
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 79 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 80 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 81 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 82 nsew signal tristate
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 83 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 84 nsew signal tristate
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 85 nsew signal tristate
flabel metal2 s 59450 0 59506 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 86 nsew signal tristate
flabel metal2 s 61106 0 61162 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 87 nsew signal tristate
flabel metal2 s 62762 0 62818 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 88 nsew signal tristate
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 89 nsew signal tristate
flabel metal2 s 66074 0 66130 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 90 nsew signal tristate
flabel metal2 s 67730 0 67786 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 91 nsew signal tristate
flabel metal2 s 69386 0 69442 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 92 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 93 nsew signal tristate
flabel metal2 s 71042 0 71098 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 94 nsew signal tristate
flabel metal2 s 72698 0 72754 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 95 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 96 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 97 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 98 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 99 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 100 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 101 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 102 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 103 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 104 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 105 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 106 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 107 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_we_i
port 108 nsew signal input
rlabel metal4 74012 43500 74012 43500 0 vccd1
rlabel metal4 71012 43500 71012 43500 0 vssd1
rlabel metal1 21758 1904 21758 1904 0 _000_
rlabel metal1 20700 2074 20700 2074 0 _001_
rlabel metal1 31648 3502 31648 3502 0 _002_
rlabel metal2 32246 4624 32246 4624 0 _003_
rlabel metal2 32890 4896 32890 4896 0 _004_
rlabel metal2 33350 4284 33350 4284 0 _005_
rlabel metal2 34914 4556 34914 4556 0 _006_
rlabel metal1 34270 4692 34270 4692 0 _007_
rlabel metal2 45954 3740 45954 3740 0 _008_
rlabel metal1 47334 3026 47334 3026 0 _009_
rlabel metal2 49082 3740 49082 3740 0 _010_
rlabel metal1 54786 5168 54786 5168 0 _011_
rlabel metal2 52946 4012 52946 4012 0 _012_
rlabel metal2 54694 4012 54694 4012 0 _013_
rlabel metal2 56258 4284 56258 4284 0 _014_
rlabel metal2 57822 4386 57822 4386 0 _015_
rlabel metal2 59478 4386 59478 4386 0 _016_
rlabel metal2 61226 4284 61226 4284 0 _017_
rlabel metal2 63250 4267 63250 4267 0 _018_
rlabel metal2 64814 4284 64814 4284 0 _019_
rlabel metal2 66470 4284 66470 4284 0 _020_
rlabel metal2 68126 4284 68126 4284 0 _021_
rlabel metal2 69874 4012 69874 4012 0 _022_
rlabel metal2 71438 4012 71438 4012 0 _023_
rlabel metal1 73094 3026 73094 3026 0 _024_
rlabel metal1 17526 2482 17526 2482 0 _025_
rlabel metal1 28014 3706 28014 3706 0 _026_
rlabel metal2 24886 4182 24886 4182 0 _027_
rlabel metal1 72588 5202 72588 5202 0 _028_
rlabel metal1 28198 2550 28198 2550 0 _029_
rlabel metal1 26404 3026 26404 3026 0 _030_
rlabel metal1 26726 3060 26726 3060 0 _031_
rlabel metal1 28428 3502 28428 3502 0 _032_
rlabel metal2 28566 4012 28566 4012 0 _033_
rlabel metal1 28106 2482 28106 2482 0 _034_
rlabel metal1 29256 1326 29256 1326 0 _035_
rlabel metal2 30038 3910 30038 3910 0 _036_
rlabel metal1 29716 3026 29716 3026 0 _037_
rlabel metal2 34730 4284 34730 4284 0 _038_
rlabel metal2 31234 4386 31234 4386 0 _039_
rlabel metal3 67091 33252 67091 33252 0 clknet_0_wb_clk_i
rlabel metal1 20010 1972 20010 1972 0 clknet_1_0__leaf_wb_clk_i
rlabel metal1 63250 53280 63250 53280 0 clknet_1_1__leaf_wb_clk_i
rlabel metal1 21068 3026 21068 3026 0 net1
rlabel metal1 43194 2312 43194 2312 0 net10
rlabel metal2 65182 1530 65182 1530 0 net100
rlabel metal1 63250 72262 63250 72262 0 net101
rlabel metal1 25852 3162 25852 3162 0 net102
rlabel metal1 63250 36405 63250 36405 0 net103
rlabel metal1 22816 1530 22816 1530 0 net104
rlabel metal1 63250 38699 63250 38699 0 net105
rlabel metal1 66700 1938 66700 1938 0 net106
rlabel metal1 63250 74590 63250 74590 0 net107
rlabel metal1 38226 1938 38226 1938 0 net108
rlabel metal1 63250 21159 63250 21159 0 net109
rlabel metal3 67091 23596 67091 23596 0 net11
rlabel metal2 67298 2244 67298 2244 0 net110
rlabel metal1 63250 76618 63250 76618 0 net111
rlabel metal1 44850 2414 44850 2414 0 net112
rlabel metal1 63250 12563 63250 12563 0 net113
rlabel metal2 20286 3910 20286 3910 0 net114
rlabel metal1 63395 40838 63395 40838 0 net115
rlabel metal1 18722 3502 18722 3502 0 net116
rlabel metal1 63395 43018 63395 43018 0 net117
rlabel metal2 69414 2108 69414 2108 0 net118
rlabel metal1 63250 78796 63250 78796 0 net119
rlabel metal3 66585 22372 66585 22372 0 net12
rlabel metal1 36754 2074 36754 2074 0 net120
rlabel metal1 63250 23337 63250 23337 0 net121
rlabel metal1 43378 1326 43378 1326 0 net122
rlabel metal1 63250 14625 63250 14625 0 net123
rlabel metal1 71668 1938 71668 1938 0 net124
rlabel metal1 63250 81008 63250 81008 0 net125
rlabel metal1 34592 3026 34592 3026 0 net126
rlabel metal1 63250 25515 63250 25515 0 net127
rlabel metal1 73140 1326 73140 1326 0 net128
rlabel metal1 63250 83186 63250 83186 0 net129
rlabel metal3 66401 23460 66401 23460 0 net13
rlabel metal1 41768 1938 41768 1938 0 net130
rlabel metal1 63250 16735 63250 16735 0 net131
rlabel metal1 33074 3026 33074 3026 0 net132
rlabel metal1 63434 25908 63434 25908 0 net133
rlabel metal1 31648 3026 31648 3026 0 net134
rlabel metal3 63687 16524 63687 16524 0 net135
rlabel metal1 29624 1938 29624 1938 0 net136
rlabel metal1 63526 26010 63526 26010 0 net137
rlabel metal1 54096 3026 54096 3026 0 net138
rlabel metal1 63250 57050 63250 57050 0 net139
rlabel metal2 20930 3332 20930 3332 0 net14
rlabel metal1 51934 1938 51934 1938 0 net140
rlabel metal1 63250 54838 63250 54838 0 net141
rlabel metal1 50186 1938 50186 1938 0 net142
rlabel metal1 63250 52694 63250 52694 0 net143
rlabel metal1 48116 1530 48116 1530 0 net144
rlabel metal1 63250 50482 63250 50482 0 net145
rlabel metal2 55062 2210 55062 2210 0 net146
rlabel metal1 63250 59194 63250 59194 0 net147
rlabel metal2 56718 1836 56718 1836 0 net148
rlabel metal1 63250 61372 63250 61372 0 net149
rlabel metal1 19458 3604 19458 3604 0 net15
rlabel metal1 59938 1938 59938 1938 0 net150
rlabel metal1 63250 65728 63250 65728 0 net151
rlabel metal1 58558 1938 58558 1938 0 net152
rlabel metal1 63250 63584 63250 63584 0 net153
rlabel metal1 35236 2414 35236 2414 0 net154
rlabel metal1 63250 44445 63250 44445 0 net155
rlabel metal1 61456 1530 61456 1530 0 net156
rlabel metal1 63250 67906 63250 67906 0 net157
rlabel metal1 27922 3162 27922 3162 0 net158
rlabel metal1 63250 34125 63250 34125 0 net159
rlabel metal1 43562 1870 43562 1870 0 net16
rlabel metal2 63618 2210 63618 2210 0 net160
rlabel metal1 63250 70084 63250 70084 0 net161
rlabel metal1 34178 2550 34178 2550 0 net162
rlabel metal1 63618 44526 63618 44526 0 net163
rlabel metal1 32108 2074 32108 2074 0 net164
rlabel metal1 63250 45003 63250 45003 0 net165
rlabel metal1 28934 1904 28934 1904 0 net166
rlabel metal1 63756 45254 63756 45254 0 net167
rlabel metal1 29210 2618 29210 2618 0 net168
rlabel metal1 63618 45730 63618 45730 0 net169
rlabel metal2 41722 2244 41722 2244 0 net17
rlabel metal1 26864 1734 26864 1734 0 net170
rlabel metal1 63250 45989 63250 45989 0 net171
rlabel metal2 25254 3060 25254 3060 0 net172
rlabel metal1 63664 43826 63664 43826 0 net173
rlabel metal1 19734 1292 19734 1292 0 net174
rlabel metal1 64032 47022 64032 47022 0 net175
rlabel metal2 20562 3332 20562 3332 0 net176
rlabel metal1 63158 47445 63158 47445 0 net177
rlabel metal1 18216 2618 18216 2618 0 net178
rlabel via3 63917 47668 63917 47668 0 net179
rlabel metal1 42136 1734 42136 1734 0 net18
rlabel metal1 22310 1938 22310 1938 0 net180
rlabel metal1 63250 22271 63250 22271 0 net181
rlabel metal1 21574 2618 21574 2618 0 net182
rlabel metal2 19826 2074 19826 2074 0 net183
rlabel metal1 63250 41873 63250 41873 0 net184
rlabel metal1 19090 2618 19090 2618 0 net185
rlabel metal1 24702 1938 24702 1938 0 net186
rlabel metal1 63250 62268 63250 62268 0 net187
rlabel metal1 24104 2618 24104 2618 0 net188
rlabel metal1 26818 1938 26818 1938 0 net189
rlabel metal1 51934 1768 51934 1768 0 net19
rlabel metal1 63250 81904 63250 81904 0 net190
rlabel metal1 25668 1530 25668 1530 0 net191
rlabel metal1 44666 1326 44666 1326 0 net192
rlabel metal1 44896 1938 44896 1938 0 net193
rlabel metal1 34960 2822 34960 2822 0 net194
rlabel metal2 33994 4250 33994 4250 0 net195
rlabel metal1 17986 1326 17986 1326 0 net196
rlabel metal2 46230 2142 46230 2142 0 net197
rlabel metal1 46000 1530 46000 1530 0 net198
rlabel metal1 44390 1360 44390 1360 0 net199
rlabel metal2 17894 3536 17894 3536 0 net2
rlabel metal1 46690 2312 46690 2312 0 net20
rlabel metal1 41216 1530 41216 1530 0 net200
rlabel metal1 39836 1870 39836 1870 0 net201
rlabel metal1 37766 1530 37766 1530 0 net202
rlabel metal1 35880 1258 35880 1258 0 net203
rlabel metal1 33948 1870 33948 1870 0 net204
rlabel metal2 32522 2244 32522 2244 0 net205
rlabel metal1 30728 1530 30728 1530 0 net206
rlabel metal1 54004 1326 54004 1326 0 net207
rlabel metal1 51428 1530 51428 1530 0 net208
rlabel metal2 29118 2108 29118 2108 0 net209
rlabel metal1 47610 2074 47610 2074 0 net21
rlabel metal2 49542 2108 49542 2108 0 net210
rlabel metal1 49496 1326 49496 1326 0 net211
rlabel metal1 54648 1938 54648 1938 0 net212
rlabel metal2 25346 2788 25346 2788 0 net213
rlabel metal2 59386 1598 59386 1598 0 net214
rlabel metal2 57270 1530 57270 1530 0 net215
rlabel metal1 64170 1530 64170 1530 0 net216
rlabel metal2 57914 2108 57914 2108 0 net217
rlabel metal2 27554 2788 27554 2788 0 net218
rlabel metal2 62422 1530 62422 1530 0 net219
rlabel metal1 66838 26350 66838 26350 0 net22
rlabel metal1 22310 1326 22310 1326 0 net220
rlabel metal2 62974 2108 62974 2108 0 net221
rlabel metal2 66102 2108 66102 2108 0 net222
rlabel metal1 68034 1870 68034 1870 0 net223
rlabel metal1 20424 2618 20424 2618 0 net224
rlabel metal1 18032 1938 18032 1938 0 net225
rlabel metal1 70104 1530 70104 1530 0 net226
rlabel metal2 71070 2108 71070 2108 0 net227
rlabel metal1 73416 1870 73416 1870 0 net228
rlabel metal1 35972 2414 35972 2414 0 net229
rlabel metal1 67114 22202 67114 22202 0 net23
rlabel metal1 33304 1190 33304 1190 0 net230
rlabel metal2 31326 2108 31326 2108 0 net231
rlabel metal2 30958 2652 30958 2652 0 net232
rlabel metal1 28244 1530 28244 1530 0 net233
rlabel metal2 26174 2176 26174 2176 0 net234
rlabel metal1 24380 2074 24380 2074 0 net235
rlabel metal2 23138 3196 23138 3196 0 net236
rlabel metal2 19918 2788 19918 2788 0 net237
rlabel metal1 17526 2074 17526 2074 0 net238
rlabel metal1 61134 2380 61134 2380 0 net24
rlabel metal1 66654 29614 66654 29614 0 net25
rlabel metal1 27738 4080 27738 4080 0 net26
rlabel metal2 66608 26860 66608 26860 0 net27
rlabel metal1 63526 2278 63526 2278 0 net28
rlabel metal2 66516 26220 66516 26220 0 net29
rlabel metal2 46046 1530 46046 1530 0 net3
rlabel metal1 66516 33422 66516 33422 0 net30
rlabel metal1 63250 2482 63250 2482 0 net31
rlabel metal1 64722 2550 64722 2550 0 net32
rlabel metal1 65826 1224 65826 1224 0 net33
rlabel metal1 66976 2006 66976 2006 0 net34
rlabel metal1 66884 39406 66884 39406 0 net35
rlabel metal1 69184 2006 69184 2006 0 net36
rlabel metal1 36570 2312 36570 2312 0 net37
rlabel metal1 71070 2006 71070 2006 0 net38
rlabel metal1 71438 1258 71438 1258 0 net39
rlabel metal1 45402 1496 45402 1496 0 net4
rlabel metal2 44666 4352 44666 4352 0 net40
rlabel metal1 27830 3400 27830 3400 0 net41
rlabel metal1 29532 3162 29532 3162 0 net42
rlabel metal2 32614 3672 32614 3672 0 net43
rlabel metal1 32936 2822 32936 2822 0 net44
rlabel metal1 34086 2822 34086 2822 0 net45
rlabel metal1 36064 3026 36064 3026 0 net46
rlabel metal1 21551 1394 21551 1394 0 net47
rlabel metal2 43010 4964 43010 4964 0 net48
rlabel metal1 68264 26962 68264 26962 0 net49
rlabel metal2 32338 4250 32338 4250 0 net5
rlabel metal1 64860 2040 64860 2040 0 net50
rlabel metal1 21252 2958 21252 2958 0 net51
rlabel metal1 20378 4148 20378 4148 0 net52
rlabel metal2 5106 1156 5106 1156 0 net53
rlabel metal2 17802 1802 17802 1802 0 net54
rlabel metal2 21482 1870 21482 1870 0 net55
rlabel metal1 37766 1326 37766 1326 0 net56
rlabel metal1 36110 3366 36110 3366 0 net57
rlabel metal2 42458 2210 42458 2210 0 net58
rlabel metal1 34270 3162 34270 3162 0 net59
rlabel metal2 19458 1054 19458 1054 0 net6
rlabel metal2 44896 1734 44896 1734 0 net60
rlabel metal1 47472 1326 47472 1326 0 net61
rlabel metal1 47794 1938 47794 1938 0 net62
rlabel metal1 48898 2890 48898 2890 0 net63
rlabel metal2 52670 2074 52670 2074 0 net64
rlabel metal2 53130 2380 53130 2380 0 net65
rlabel metal1 22862 2448 22862 2448 0 net66
rlabel metal1 55062 2822 55062 2822 0 net67
rlabel metal2 56442 2380 56442 2380 0 net68
rlabel metal2 58006 2074 58006 2074 0 net69
rlabel metal2 24978 4828 24978 4828 0 net7
rlabel metal1 60030 2822 60030 2822 0 net70
rlabel metal2 61410 2380 61410 2380 0 net71
rlabel metal2 63066 2074 63066 2074 0 net72
rlabel metal2 64630 2380 64630 2380 0 net73
rlabel metal2 66286 2074 66286 2074 0 net74
rlabel metal2 68310 2074 68310 2074 0 net75
rlabel metal2 69690 2380 69690 2380 0 net76
rlabel metal1 24150 1258 24150 1258 0 net77
rlabel metal2 71254 2074 71254 2074 0 net78
rlabel metal2 73278 2074 73278 2074 0 net79
rlabel metal2 27094 4590 27094 4590 0 net8
rlabel metal1 26726 1258 26726 1258 0 net80
rlabel metal1 27968 1326 27968 1326 0 net81
rlabel metal1 29762 1972 29762 1972 0 net82
rlabel metal1 30498 1292 30498 1292 0 net83
rlabel metal1 32522 3128 32522 3128 0 net84
rlabel metal1 33442 2958 33442 2958 0 net85
rlabel metal2 35650 1156 35650 1156 0 net86
rlabel metal1 63618 49631 63618 49631 0 net87
rlabel metal1 63250 43713 63250 43713 0 net88
rlabel metal1 63250 42543 63250 42543 0 net89
rlabel metal2 28934 4726 28934 4726 0 net9
rlabel metal1 63250 50114 63250 50114 0 net90
rlabel metal1 63441 52094 63441 52094 0 net91
rlabel metal1 63250 52289 63250 52289 0 net92
rlabel metal1 63441 48715 63441 48715 0 net93
rlabel metal1 66424 47022 66424 47022 0 net94
rlabel metal1 66378 46954 66378 46954 0 net95
rlabel metal2 39146 2210 39146 2210 0 net96
rlabel metal1 63250 18981 63250 18981 0 net97
rlabel metal1 46920 1938 46920 1938 0 net98
rlabel metal1 55752 5542 55752 5542 0 net99
rlabel metal1 63250 43283 63250 43283 0 ram_controller.DO\[0\]
rlabel metal1 63441 21470 63441 21470 0 ram_controller.DO\[10\]
rlabel metal1 63250 19209 63250 19209 0 ram_controller.DO\[11\]
rlabel metal1 63250 17031 63250 17031 0 ram_controller.DO\[12\]
rlabel metal1 63250 14853 63250 14853 0 ram_controller.DO\[13\]
rlabel via2 64906 12733 64906 12733 0 ram_controller.DO\[14\]
rlabel metal2 27554 5882 27554 5882 0 ram_controller.DO\[15\]
rlabel metal1 63250 50288 63250 50288 0 ram_controller.DO\[16\]
rlabel metal1 63158 52548 63158 52548 0 ram_controller.DO\[17\]
rlabel metal1 63158 54644 63158 54644 0 ram_controller.DO\[18\]
rlabel metal1 63250 56754 63250 56754 0 ram_controller.DO\[19\]
rlabel metal1 63250 41023 63250 41023 0 ram_controller.DO\[1\]
rlabel metal1 63250 59048 63250 59048 0 ram_controller.DO\[20\]
rlabel metal1 63618 25908 63618 25908 0 ram_controller.DO\[21\]
rlabel metal1 63250 63404 63250 63404 0 ram_controller.DO\[22\]
rlabel metal1 63250 65466 63250 65466 0 ram_controller.DO\[23\]
rlabel metal1 63250 67678 63250 67678 0 ram_controller.DO\[24\]
rlabel metal3 63457 26180 63457 26180 0 ram_controller.DO\[25\]
rlabel metal1 63250 72000 63250 72000 0 ram_controller.DO\[26\]
rlabel metal1 63250 74178 63250 74178 0 ram_controller.DO\[27\]
rlabel metal1 63250 76472 63250 76472 0 ram_controller.DO\[28\]
rlabel metal1 63250 78636 63250 78636 0 ram_controller.DO\[29\]
rlabel metal1 63441 38910 63441 38910 0 ram_controller.DO\[2\]
rlabel metal1 63250 80814 63250 80814 0 ram_controller.DO\[30\]
rlabel metal1 63250 82992 63250 82992 0 ram_controller.DO\[31\]
rlabel metal1 63250 36633 63250 36633 0 ram_controller.DO\[3\]
rlabel metal1 63250 34571 63250 34571 0 ram_controller.DO\[4\]
rlabel metal1 63250 32277 63250 32277 0 ram_controller.DO\[5\]
rlabel metal1 63250 30099 63250 30099 0 ram_controller.DO\[6\]
rlabel metal1 63250 27921 63250 27921 0 ram_controller.DO\[7\]
rlabel metal1 63250 25743 63250 25743 0 ram_controller.DO\[8\]
rlabel metal1 63250 23565 63250 23565 0 ram_controller.DO\[9\]
rlabel metal3 63227 48756 63227 48756 0 ram_controller.EN
rlabel metal3 64009 48076 64009 48076 0 ram_controller.R_WB
rlabel metal2 20654 3196 20654 3196 0 ram_controller.wbs_ack_o
rlabel metal2 3174 1010 3174 1010 0 sram_selected
rlabel metal2 14766 2047 14766 2047 0 wb_clk_i
rlabel metal2 15318 1044 15318 1044 0 wb_rst_i
rlabel metal2 15870 1010 15870 1010 0 wbs_ack_o
rlabel metal2 18078 1316 18078 1316 0 wbs_adr_i[0]
rlabel metal2 43470 1588 43470 1588 0 wbs_adr_i[14]
rlabel metal2 45126 1010 45126 1010 0 wbs_adr_i[15]
rlabel metal2 20286 1010 20286 1010 0 wbs_adr_i[1]
rlabel metal1 22540 3502 22540 3502 0 wbs_adr_i[2]
rlabel metal2 24702 1316 24702 1316 0 wbs_adr_i[3]
rlabel metal2 26910 1588 26910 1588 0 wbs_adr_i[4]
rlabel metal2 28566 840 28566 840 0 wbs_adr_i[5]
rlabel metal1 30268 2958 30268 2958 0 wbs_adr_i[6]
rlabel metal2 31878 823 31878 823 0 wbs_adr_i[7]
rlabel metal2 33534 1044 33534 1044 0 wbs_adr_i[8]
rlabel metal2 35190 823 35190 823 0 wbs_adr_i[9]
rlabel metal2 16422 1350 16422 1350 0 wbs_cyc_i
rlabel metal1 18860 2958 18860 2958 0 wbs_dat_i[0]
rlabel metal2 37398 1044 37398 1044 0 wbs_dat_i[10]
rlabel metal2 39054 1350 39054 1350 0 wbs_dat_i[11]
rlabel metal2 40710 823 40710 823 0 wbs_dat_i[12]
rlabel metal2 42366 1588 42366 1588 0 wbs_dat_i[13]
rlabel metal2 44022 1010 44022 1010 0 wbs_dat_i[14]
rlabel metal2 45678 1350 45678 1350 0 wbs_dat_i[15]
rlabel metal2 47334 1588 47334 1588 0 wbs_dat_i[16]
rlabel metal2 48990 1010 48990 1010 0 wbs_dat_i[17]
rlabel metal2 50646 1044 50646 1044 0 wbs_dat_i[18]
rlabel metal2 52302 976 52302 976 0 wbs_dat_i[19]
rlabel metal2 20838 1622 20838 1622 0 wbs_dat_i[1]
rlabel metal2 53958 1588 53958 1588 0 wbs_dat_i[20]
rlabel metal2 55614 1316 55614 1316 0 wbs_dat_i[21]
rlabel metal2 57270 959 57270 959 0 wbs_dat_i[22]
rlabel metal2 58926 1010 58926 1010 0 wbs_dat_i[23]
rlabel metal2 60582 1316 60582 1316 0 wbs_dat_i[24]
rlabel metal2 62238 1027 62238 1027 0 wbs_dat_i[25]
rlabel metal2 63894 1044 63894 1044 0 wbs_dat_i[26]
rlabel metal2 65550 1588 65550 1588 0 wbs_dat_i[27]
rlabel metal2 67206 1350 67206 1350 0 wbs_dat_i[28]
rlabel metal2 68862 1044 68862 1044 0 wbs_dat_i[29]
rlabel metal1 23414 2958 23414 2958 0 wbs_dat_i[2]
rlabel metal2 70518 1588 70518 1588 0 wbs_dat_i[30]
rlabel metal2 72174 823 72174 823 0 wbs_dat_i[31]
rlabel metal2 25254 1588 25254 1588 0 wbs_dat_i[3]
rlabel metal2 27462 1588 27462 1588 0 wbs_dat_i[4]
rlabel metal2 29118 1027 29118 1027 0 wbs_dat_i[5]
rlabel metal2 30774 823 30774 823 0 wbs_dat_i[6]
rlabel metal2 32430 1316 32430 1316 0 wbs_dat_i[7]
rlabel metal2 34086 1350 34086 1350 0 wbs_dat_i[8]
rlabel metal2 35742 976 35742 976 0 wbs_dat_i[9]
rlabel metal2 19182 1078 19182 1078 0 wbs_dat_o[0]
rlabel metal2 37950 1078 37950 1078 0 wbs_dat_o[10]
rlabel metal2 39606 1010 39606 1010 0 wbs_dat_o[11]
rlabel metal2 41262 1078 41262 1078 0 wbs_dat_o[12]
rlabel metal2 42918 874 42918 874 0 wbs_dat_o[13]
rlabel metal2 44574 823 44574 823 0 wbs_dat_o[14]
rlabel metal2 46230 1078 46230 1078 0 wbs_dat_o[15]
rlabel metal2 47886 1316 47886 1316 0 wbs_dat_o[16]
rlabel metal2 49542 823 49542 823 0 wbs_dat_o[17]
rlabel metal2 51198 1010 51198 1010 0 wbs_dat_o[18]
rlabel metal2 52854 1316 52854 1316 0 wbs_dat_o[19]
rlabel metal2 21390 1588 21390 1588 0 wbs_dat_o[1]
rlabel metal2 54510 823 54510 823 0 wbs_dat_o[20]
rlabel metal2 56166 1316 56166 1316 0 wbs_dat_o[21]
rlabel metal2 57822 1010 57822 1010 0 wbs_dat_o[22]
rlabel metal2 59478 1078 59478 1078 0 wbs_dat_o[23]
rlabel metal2 61134 1316 61134 1316 0 wbs_dat_o[24]
rlabel metal2 62790 1078 62790 1078 0 wbs_dat_o[25]
rlabel metal2 64446 823 64446 823 0 wbs_dat_o[26]
rlabel metal2 66102 1010 66102 1010 0 wbs_dat_o[27]
rlabel metal2 67758 1078 67758 1078 0 wbs_dat_o[28]
rlabel metal2 69414 1282 69414 1282 0 wbs_dat_o[29]
rlabel metal2 23598 1010 23598 1010 0 wbs_dat_o[2]
rlabel metal2 71070 1078 71070 1078 0 wbs_dat_o[30]
rlabel metal2 72726 976 72726 976 0 wbs_dat_o[31]
rlabel metal2 25806 1010 25806 1010 0 wbs_dat_o[3]
rlabel metal2 28014 1078 28014 1078 0 wbs_dat_o[4]
rlabel metal2 29670 823 29670 823 0 wbs_dat_o[5]
rlabel metal2 31326 1010 31326 1010 0 wbs_dat_o[6]
rlabel metal2 32982 1010 32982 1010 0 wbs_dat_o[7]
rlabel metal2 34638 1316 34638 1316 0 wbs_dat_o[8]
rlabel metal2 36294 1010 36294 1010 0 wbs_dat_o[9]
rlabel metal2 19734 1622 19734 1622 0 wbs_sel_i[0]
rlabel metal2 21942 823 21942 823 0 wbs_sel_i[1]
rlabel metal2 24150 823 24150 823 0 wbs_sel_i[2]
rlabel metal2 26358 1044 26358 1044 0 wbs_sel_i[3]
rlabel metal2 16974 1588 16974 1588 0 wbs_stb_i
rlabel metal2 17526 1044 17526 1044 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 76000 87000
<< end >>
