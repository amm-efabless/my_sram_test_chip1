magic
tech sky130A
magscale 1 2
timestamp 1715271074
<< viali >>
rect 65625 52445 65659 52479
rect 65901 52445 65935 52479
rect 65625 50269 65659 50303
rect 65625 49589 65659 49623
rect 65625 49181 65659 49215
rect 65625 47005 65659 47039
rect 65901 46937 65935 46971
rect 65625 43741 65659 43775
rect 68017 42721 68051 42755
rect 65625 42653 65659 42687
rect 68661 42653 68695 42687
rect 67097 41769 67131 41803
rect 67741 41565 67775 41599
rect 66453 40681 66487 40715
rect 67097 40477 67131 40511
rect 65625 39593 65659 39627
rect 66269 39389 66303 39423
rect 65625 38505 65659 38539
rect 66269 38301 66303 38335
rect 66269 37213 66303 37247
rect 65625 37145 65659 37179
rect 65625 36329 65659 36363
rect 66269 36125 66303 36159
rect 66545 35717 66579 35751
rect 65809 35649 65843 35683
rect 65625 35241 65659 35275
rect 66269 35037 66303 35071
rect 66913 34153 66947 34187
rect 65625 33881 65659 33915
rect 65625 33609 65659 33643
rect 66269 33405 66303 33439
rect 65625 33065 65659 33099
rect 66269 32861 66303 32895
rect 65625 31977 65659 32011
rect 66269 31773 66303 31807
rect 65625 30889 65659 30923
rect 66269 30685 66303 30719
rect 65625 29801 65659 29835
rect 66269 29597 66303 29631
rect 65625 28713 65659 28747
rect 66269 28509 66303 28543
rect 65625 27557 65659 27591
rect 66269 27421 66303 27455
rect 65809 26945 65843 26979
rect 66361 26877 66395 26911
rect 65625 26537 65659 26571
rect 66269 26333 66303 26367
rect 65625 24361 65659 24395
rect 66269 24157 66303 24191
rect 65625 23817 65659 23851
rect 66269 23613 66303 23647
rect 65625 23273 65659 23307
rect 66269 23069 66303 23103
rect 23673 5865 23707 5899
rect 24133 5865 24167 5899
rect 49617 5865 49651 5899
rect 51089 5865 51123 5899
rect 56149 5797 56183 5831
rect 23305 5729 23339 5763
rect 23765 5729 23799 5763
rect 24317 5729 24351 5763
rect 24685 5729 24719 5763
rect 48237 5729 48271 5763
rect 48881 5729 48915 5763
rect 48973 5729 49007 5763
rect 54769 5729 54803 5763
rect 56517 5729 56551 5763
rect 57805 5729 57839 5763
rect 58173 5729 58207 5763
rect 59737 5729 59771 5763
rect 61669 5729 61703 5763
rect 62957 5729 62991 5763
rect 65073 5729 65107 5763
rect 66177 5729 66211 5763
rect 68477 5729 68511 5763
rect 23489 5661 23523 5695
rect 23949 5661 23983 5695
rect 24501 5661 24535 5695
rect 24777 5661 24811 5695
rect 24961 5661 24995 5695
rect 25881 5661 25915 5695
rect 25973 5661 26007 5695
rect 26157 5661 26191 5695
rect 40417 5661 40451 5695
rect 42349 5661 42383 5695
rect 43821 5661 43855 5695
rect 44465 5661 44499 5695
rect 44925 5661 44959 5695
rect 45661 5661 45695 5695
rect 46305 5661 46339 5695
rect 46397 5661 46431 5695
rect 47041 5661 47075 5695
rect 47501 5661 47535 5695
rect 50445 5661 50479 5695
rect 51273 5661 51307 5695
rect 51917 5661 51951 5695
rect 52653 5661 52687 5695
rect 53389 5661 53423 5695
rect 54033 5661 54067 5695
rect 54217 5661 54251 5695
rect 55321 5661 55355 5695
rect 55873 5661 55907 5695
rect 56333 5661 56367 5695
rect 57989 5661 58023 5695
rect 59553 5661 59587 5695
rect 61485 5661 61519 5695
rect 63141 5661 63175 5695
rect 64889 5661 64923 5695
rect 66361 5661 66395 5695
rect 68293 5661 68327 5695
rect 37013 5593 37047 5627
rect 43545 5593 43579 5627
rect 25145 5525 25179 5559
rect 35725 5525 35759 5559
rect 41705 5525 41739 5559
rect 45569 5525 45603 5559
rect 48145 5525 48179 5559
rect 53297 5525 53331 5559
rect 59369 5525 59403 5559
rect 61301 5525 61335 5559
rect 63325 5525 63359 5559
rect 64705 5525 64739 5559
rect 66545 5525 66579 5559
rect 68109 5525 68143 5559
rect 27905 5321 27939 5355
rect 41061 5321 41095 5355
rect 24409 5185 24443 5219
rect 24869 5185 24903 5219
rect 25605 5185 25639 5219
rect 26065 5185 26099 5219
rect 26525 5185 26559 5219
rect 27261 5185 27295 5219
rect 27721 5185 27755 5219
rect 28273 5185 28307 5219
rect 28917 5185 28951 5219
rect 29561 5185 29595 5219
rect 30113 5185 30147 5219
rect 30297 5185 30331 5219
rect 30665 5185 30699 5219
rect 30849 5185 30883 5219
rect 42993 5185 43027 5219
rect 44189 5185 44223 5219
rect 46213 5185 46247 5219
rect 46305 5185 46339 5219
rect 47225 5185 47259 5219
rect 53113 5185 53147 5219
rect 54769 5185 54803 5219
rect 54861 5185 54895 5219
rect 70225 5185 70259 5219
rect 71697 5185 71731 5219
rect 73445 5185 73479 5219
rect 73537 5185 73571 5219
rect 24225 5117 24259 5151
rect 25421 5117 25455 5151
rect 25881 5117 25915 5151
rect 26341 5117 26375 5151
rect 27077 5117 27111 5151
rect 27537 5117 27571 5151
rect 28457 5117 28491 5151
rect 29101 5117 29135 5151
rect 29745 5117 29779 5151
rect 40417 5117 40451 5151
rect 41521 5117 41555 5151
rect 42165 5117 42199 5151
rect 44557 5117 44591 5151
rect 45385 5117 45419 5151
rect 46581 5117 46615 5151
rect 47501 5117 47535 5151
rect 48145 5117 48179 5151
rect 49157 5117 49191 5151
rect 49801 5117 49835 5151
rect 53297 5117 53331 5151
rect 70409 5117 70443 5151
rect 71881 5117 71915 5151
rect 24685 5049 24719 5083
rect 25789 5049 25823 5083
rect 27445 5049 27479 5083
rect 45109 5049 45143 5083
rect 24593 4981 24627 5015
rect 26249 4981 26283 5015
rect 26709 4981 26743 5015
rect 28089 4981 28123 5015
rect 28733 4981 28767 5015
rect 29377 4981 29411 5015
rect 29929 4981 29963 5015
rect 30481 4981 30515 5015
rect 46029 4981 46063 5015
rect 46489 4981 46523 5015
rect 52929 4981 52963 5015
rect 54585 4981 54619 5015
rect 70041 4981 70075 5015
rect 71513 4981 71547 5015
rect 73261 4981 73295 5015
rect 61117 4777 61151 4811
rect 44097 4641 44131 4675
rect 33977 4573 34011 4607
rect 34253 4573 34287 4607
rect 41245 4573 41279 4607
rect 41981 4573 42015 4607
rect 43453 4573 43487 4607
rect 44281 4573 44315 4607
rect 46765 4573 46799 4607
rect 46857 4573 46891 4607
rect 61209 4573 61243 4607
rect 41889 4437 41923 4471
rect 42625 4437 42659 4471
rect 44005 4437 44039 4471
rect 44465 4437 44499 4471
rect 47041 4437 47075 4471
rect 19717 4097 19751 4131
rect 27629 4097 27663 4131
rect 30849 4097 30883 4131
rect 31309 4097 31343 4131
rect 34713 4097 34747 4131
rect 34897 4097 34931 4131
rect 19533 4029 19567 4063
rect 29745 4029 29779 4063
rect 27721 3893 27755 3927
rect 30389 3893 30423 3927
rect 20269 3689 20303 3723
rect 26065 3689 26099 3723
rect 26249 3689 26283 3723
rect 31401 3689 31435 3723
rect 32413 3689 32447 3723
rect 19441 3553 19475 3587
rect 23673 3553 23707 3587
rect 24961 3553 24995 3587
rect 25605 3553 25639 3587
rect 19165 3485 19199 3519
rect 20177 3485 20211 3519
rect 20821 3485 20855 3519
rect 22569 3485 22603 3519
rect 23489 3485 23523 3519
rect 25237 3485 25271 3519
rect 25789 3485 25823 3519
rect 28089 3485 28123 3519
rect 31217 3485 31251 3519
rect 31677 3485 31711 3519
rect 32229 3485 32263 3519
rect 32873 3485 32907 3519
rect 19901 3417 19935 3451
rect 25881 3417 25915 3451
rect 26097 3417 26131 3451
rect 27721 3417 27755 3451
rect 23213 3349 23247 3383
rect 23305 3349 23339 3383
rect 27629 3349 27663 3383
rect 27905 3349 27939 3383
rect 31861 3349 31895 3383
rect 33057 3349 33091 3383
rect 20545 3145 20579 3179
rect 20913 3145 20947 3179
rect 21281 3145 21315 3179
rect 25881 3145 25915 3179
rect 28089 3145 28123 3179
rect 29469 3145 29503 3179
rect 30205 3145 30239 3179
rect 31493 3145 31527 3179
rect 33517 3145 33551 3179
rect 37013 3145 37047 3179
rect 17877 3077 17911 3111
rect 21122 3077 21156 3111
rect 35909 3077 35943 3111
rect 54585 3077 54619 3111
rect 18153 3009 18187 3043
rect 20637 3009 20671 3043
rect 21373 3009 21407 3043
rect 23121 3009 23155 3043
rect 26157 3009 26191 3043
rect 26709 3009 26743 3043
rect 26893 3009 26927 3043
rect 28549 3009 28583 3043
rect 29101 3009 29135 3043
rect 29561 3009 29595 3043
rect 29745 3009 29779 3043
rect 30021 3009 30055 3043
rect 31585 3009 31619 3043
rect 32045 3009 32079 3043
rect 32597 3009 32631 3043
rect 32965 3009 32999 3043
rect 33333 3009 33367 3043
rect 33793 3009 33827 3043
rect 34069 3009 34103 3043
rect 34529 3009 34563 3043
rect 34897 3009 34931 3043
rect 35725 3009 35759 3043
rect 36277 3009 36311 3043
rect 36829 3009 36863 3043
rect 45937 3009 45971 3043
rect 47501 3009 47535 3043
rect 49065 3009 49099 3043
rect 52929 3009 52963 3043
rect 54217 3009 54251 3043
rect 54677 3009 54711 3043
rect 56241 3009 56275 3043
rect 57805 3009 57839 3043
rect 59461 3009 59495 3043
rect 61209 3009 61243 3043
rect 63233 3009 63267 3043
rect 64797 3009 64831 3043
rect 66453 3009 66487 3043
rect 68109 3009 68143 3043
rect 69857 3009 69891 3043
rect 71421 3009 71455 3043
rect 72893 3009 72927 3043
rect 18981 2941 19015 2975
rect 19165 2941 19199 2975
rect 19901 2941 19935 2975
rect 21005 2941 21039 2975
rect 21741 2941 21775 2975
rect 23765 2941 23799 2975
rect 24317 2941 24351 2975
rect 25329 2941 25363 2975
rect 27077 2941 27111 2975
rect 27537 2941 27571 2975
rect 28825 2941 28859 2975
rect 30297 2941 30331 2975
rect 30941 2941 30975 2975
rect 32229 2941 32263 2975
rect 35173 2941 35207 2975
rect 22477 2873 22511 2907
rect 29929 2873 29963 2907
rect 35081 2873 35115 2907
rect 47685 2873 47719 2907
rect 18429 2805 18463 2839
rect 19809 2805 19843 2839
rect 21465 2805 21499 2839
rect 22385 2805 22419 2839
rect 23213 2805 23247 2839
rect 24961 2805 24995 2839
rect 25973 2805 26007 2839
rect 26525 2805 26559 2839
rect 28365 2805 28399 2839
rect 34253 2805 34287 2839
rect 46121 2805 46155 2839
rect 49249 2805 49283 2839
rect 53113 2805 53147 2839
rect 54861 2805 54895 2839
rect 56425 2805 56459 2839
rect 57989 2805 58023 2839
rect 59645 2805 59679 2839
rect 61393 2805 61427 2839
rect 63049 2805 63083 2839
rect 64613 2805 64647 2839
rect 66269 2805 66303 2839
rect 68293 2805 68327 2839
rect 69673 2805 69707 2839
rect 71237 2805 71271 2839
rect 73077 2805 73111 2839
rect 18245 2601 18279 2635
rect 18981 2601 19015 2635
rect 19901 2601 19935 2635
rect 19993 2601 20027 2635
rect 21373 2601 21407 2635
rect 24133 2601 24167 2635
rect 25237 2601 25271 2635
rect 25329 2601 25363 2635
rect 27537 2601 27571 2635
rect 29285 2601 29319 2635
rect 31677 2601 31711 2635
rect 33149 2601 33183 2635
rect 34253 2601 34287 2635
rect 47133 2601 47167 2635
rect 53941 2601 53975 2635
rect 56057 2601 56091 2635
rect 63325 2601 63359 2635
rect 39313 2533 39347 2567
rect 44373 2533 44407 2567
rect 18429 2465 18463 2499
rect 20637 2465 20671 2499
rect 30941 2465 30975 2499
rect 60749 2465 60783 2499
rect 67465 2465 67499 2499
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 17601 2397 17635 2431
rect 19349 2397 19383 2431
rect 20729 2397 20763 2431
rect 21649 2397 21683 2431
rect 22845 2397 22879 2431
rect 22937 2397 22971 2431
rect 23581 2397 23615 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 26065 2397 26099 2431
rect 27353 2397 27387 2431
rect 28089 2397 28123 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 30021 2397 30055 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 32505 2397 32539 2431
rect 33609 2397 33643 2431
rect 35173 2397 35207 2431
rect 35265 2397 35299 2431
rect 35909 2397 35943 2431
rect 36001 2397 36035 2431
rect 36553 2397 36587 2431
rect 42441 2397 42475 2431
rect 43729 2397 43763 2431
rect 44741 2397 44775 2431
rect 44925 2397 44959 2431
rect 45569 2397 45603 2431
rect 46213 2397 46247 2431
rect 47409 2397 47443 2431
rect 49065 2397 49099 2431
rect 53389 2397 53423 2431
rect 54125 2397 54159 2431
rect 55689 2397 55723 2431
rect 57345 2397 57379 2431
rect 62313 2397 62347 2431
rect 65625 2397 65659 2431
rect 67741 2397 67775 2431
rect 69949 2397 69983 2431
rect 70685 2397 70719 2431
rect 23213 2329 23247 2363
rect 34897 2329 34931 2363
rect 39497 2329 39531 2363
rect 43085 2329 43119 2363
rect 47225 2329 47259 2363
rect 55321 2329 55355 2363
rect 56149 2329 56183 2363
rect 61025 2329 61059 2363
rect 63417 2329 63451 2363
rect 17233 2261 17267 2295
rect 17325 2261 17359 2295
rect 26709 2261 26743 2295
rect 26801 2261 26835 2295
rect 28549 2261 28583 2295
rect 29469 2261 29503 2295
rect 30297 2261 30331 2295
rect 31769 2261 31803 2295
rect 44557 2261 44591 2295
rect 46765 2261 46799 2295
rect 48053 2261 48087 2295
rect 49709 2261 49743 2295
rect 54769 2261 54803 2295
rect 57989 2261 58023 2295
rect 62957 2261 62991 2295
rect 66269 2261 66303 2295
rect 69305 2261 69339 2295
rect 71329 2261 71363 2295
rect 16405 2057 16439 2091
rect 17417 2057 17451 2091
rect 18153 2057 18187 2091
rect 24133 2057 24167 2091
rect 25697 2057 25731 2091
rect 26709 2057 26743 2091
rect 31861 2057 31895 2091
rect 32505 2057 32539 2091
rect 34621 2057 34655 2091
rect 36829 2057 36863 2091
rect 39129 2057 39163 2091
rect 41981 2057 42015 2091
rect 44741 2057 44775 2091
rect 50537 2057 50571 2091
rect 55045 2057 55079 2091
rect 58909 2057 58943 2091
rect 63601 2057 63635 2091
rect 67281 2057 67315 2091
rect 20269 1989 20303 2023
rect 28089 1989 28123 2023
rect 67005 1989 67039 2023
rect 69121 1989 69155 2023
rect 71973 1989 72007 2023
rect 16221 1921 16255 1955
rect 17601 1921 17635 1955
rect 21465 1921 21499 1955
rect 22201 1921 22235 1955
rect 24409 1921 24443 1955
rect 25881 1921 25915 1955
rect 26157 1921 26191 1955
rect 26893 1921 26927 1955
rect 28917 1921 28951 1955
rect 29101 1921 29135 1955
rect 29653 1921 29687 1955
rect 29745 1921 29779 1955
rect 31309 1921 31343 1955
rect 33333 1921 33367 1955
rect 34805 1921 34839 1955
rect 38117 1921 38151 1955
rect 38301 1921 38335 1955
rect 40417 1921 40451 1955
rect 41705 1921 41739 1955
rect 41797 1921 41831 1955
rect 42717 1921 42751 1955
rect 42993 1921 43027 1955
rect 44741 1921 44775 1955
rect 45385 1921 45419 1955
rect 46765 1921 46799 1955
rect 46949 1921 46983 1955
rect 47961 1921 47995 1955
rect 49525 1921 49559 1955
rect 50077 1921 50111 1955
rect 50261 1921 50295 1955
rect 51825 1921 51859 1955
rect 52009 1921 52043 1955
rect 53113 1921 53147 1955
rect 54493 1921 54527 1955
rect 56425 1921 56459 1955
rect 57897 1921 57931 1955
rect 58449 1921 58483 1955
rect 58633 1921 58667 1955
rect 59829 1921 59863 1955
rect 60013 1921 60047 1955
rect 61393 1921 61427 1955
rect 62957 1921 62991 1955
rect 64613 1921 64647 1955
rect 66085 1921 66119 1955
rect 66637 1921 66671 1955
rect 66729 1921 66763 1955
rect 68661 1921 68695 1955
rect 69397 1921 69431 1955
rect 69673 1921 69707 1955
rect 71053 1921 71087 1955
rect 71605 1921 71639 1955
rect 71697 1921 71731 1955
rect 16865 1853 16899 1887
rect 18245 1853 18279 1887
rect 19717 1853 19751 1887
rect 19993 1853 20027 1887
rect 23213 1853 23247 1887
rect 23581 1853 23615 1887
rect 25421 1853 25455 1887
rect 28733 1853 28767 1887
rect 30389 1853 30423 1887
rect 33149 1853 33183 1887
rect 33885 1853 33919 1887
rect 33977 1853 34011 1887
rect 35173 1853 35207 1887
rect 36185 1853 36219 1887
rect 37565 1853 37599 1887
rect 39773 1853 39807 1887
rect 39865 1853 39899 1887
rect 41153 1853 41187 1887
rect 43453 1853 43487 1887
rect 45477 1853 45511 1887
rect 46029 1853 46063 1887
rect 46213 1853 46247 1887
rect 48421 1853 48455 1887
rect 51273 1853 51307 1887
rect 53389 1853 53423 1887
rect 55597 1853 55631 1887
rect 56701 1853 56735 1887
rect 59277 1853 59311 1887
rect 60565 1853 60599 1887
rect 61669 1853 61703 1887
rect 63877 1853 63911 1887
rect 64981 1853 65015 1887
rect 67925 1853 67959 1887
rect 68109 1853 68143 1887
rect 69949 1853 69983 1887
rect 72341 1853 72375 1887
rect 72985 1853 73019 1887
rect 73813 1853 73847 1887
rect 52285 1785 52319 1819
rect 60289 1785 60323 1819
rect 38577 1717 38611 1751
rect 42533 1717 42567 1751
rect 47133 1717 47167 1751
rect 56149 1717 56183 1751
rect 61117 1717 61151 1751
rect 64429 1717 64463 1751
rect 73261 1717 73295 1751
rect 22661 1513 22695 1547
rect 25237 1513 25271 1547
rect 27813 1513 27847 1547
rect 30389 1513 30423 1547
rect 37933 1513 37967 1547
rect 41245 1513 41279 1547
rect 46397 1513 46431 1547
rect 47133 1513 47167 1547
rect 51549 1513 51583 1547
rect 61853 1513 61887 1547
rect 64429 1513 64463 1547
rect 70225 1513 70259 1547
rect 21005 1377 21039 1411
rect 28365 1377 28399 1411
rect 38485 1377 38519 1411
rect 42809 1377 42843 1411
rect 45385 1377 45419 1411
rect 47961 1377 47995 1411
rect 50537 1377 50571 1411
rect 60841 1377 60875 1411
rect 63417 1377 63451 1411
rect 68569 1377 68603 1411
rect 71605 1377 71639 1411
rect 5089 1309 5123 1343
rect 15393 1309 15427 1343
rect 15853 1309 15887 1343
rect 17785 1309 17819 1343
rect 18061 1309 18095 1343
rect 18337 1309 18371 1343
rect 19717 1309 19751 1343
rect 19809 1309 19843 1343
rect 22017 1309 22051 1343
rect 24133 1309 24167 1343
rect 24685 1309 24719 1343
rect 26709 1309 26743 1343
rect 27261 1309 27295 1343
rect 28089 1309 28123 1343
rect 29469 1309 29503 1343
rect 29837 1309 29871 1343
rect 30481 1309 30515 1343
rect 32413 1309 32447 1343
rect 33241 1309 33275 1343
rect 34989 1309 35023 1343
rect 35633 1309 35667 1343
rect 37381 1309 37415 1343
rect 38025 1309 38059 1343
rect 39773 1309 39807 1343
rect 41797 1309 41831 1343
rect 42441 1309 42475 1343
rect 43821 1309 43855 1343
rect 44465 1309 44499 1343
rect 44557 1309 44591 1343
rect 44925 1309 44959 1343
rect 46949 1309 46983 1343
rect 47317 1309 47351 1343
rect 47501 1309 47535 1343
rect 48973 1309 49007 1343
rect 49525 1309 49559 1343
rect 50077 1309 50111 1343
rect 52101 1309 52135 1343
rect 52653 1309 52687 1343
rect 54125 1309 54159 1343
rect 54677 1309 54711 1343
rect 55229 1309 55263 1343
rect 56701 1309 56735 1343
rect 57253 1309 57287 1343
rect 57989 1309 58023 1343
rect 59369 1309 59403 1343
rect 59921 1309 59955 1343
rect 60381 1309 60415 1343
rect 62405 1309 62439 1343
rect 63049 1309 63083 1343
rect 64981 1309 65015 1343
rect 65533 1309 65567 1343
rect 66269 1309 66303 1343
rect 68293 1309 68327 1343
rect 69581 1309 69615 1343
rect 71237 1309 71271 1343
rect 73077 1309 73111 1343
rect 73261 1309 73295 1343
rect 3893 1241 3927 1275
rect 16773 1241 16807 1275
rect 19441 1241 19475 1275
rect 23213 1241 23247 1275
rect 25789 1241 25823 1275
rect 31401 1241 31435 1275
rect 33977 1241 34011 1275
rect 35541 1241 35575 1275
rect 36553 1241 36587 1275
rect 40693 1241 40727 1275
rect 53573 1241 53607 1275
rect 56149 1241 56183 1275
rect 58817 1241 58851 1275
rect 65809 1241 65843 1275
rect 67097 1241 67131 1275
rect 72801 1241 72835 1275
rect 74181 1241 74215 1275
rect 15577 1173 15611 1207
rect 16405 1173 16439 1207
rect 29653 1173 29687 1207
rect 32965 1173 32999 1207
rect 44741 1173 44775 1207
<< metal1 >>
rect 65320 85978 74980 86000
rect 65320 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74980 85978
rect 65320 85904 74980 85926
rect 65320 85434 74980 85456
rect 65320 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 74980 85434
rect 65320 85360 74980 85382
rect 65320 84890 74980 84912
rect 65320 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74980 84890
rect 65320 84816 74980 84838
rect 65320 84346 74980 84368
rect 65320 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 74980 84346
rect 65320 84272 74980 84294
rect 64874 84232 64880 84244
rect 63236 84204 64880 84232
rect 64874 84192 64880 84204
rect 64932 84192 64938 84244
rect 65320 83802 74980 83824
rect 65320 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74980 83802
rect 65320 83728 74980 83750
rect 65320 83258 74980 83280
rect 63236 83144 63264 83256
rect 65320 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 74980 83258
rect 65320 83184 74980 83206
rect 66990 83144 66996 83156
rect 63236 83116 66996 83144
rect 66990 83104 66996 83116
rect 67048 83104 67054 83156
rect 69658 83008 69664 83020
rect 63236 82980 69664 83008
rect 69658 82968 69664 82980
rect 69716 82968 69722 83020
rect 65320 82714 74980 82736
rect 65320 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74980 82714
rect 65320 82640 74980 82662
rect 65320 82170 74980 82192
rect 65320 82118 71858 82170
rect 71910 82118 71922 82170
rect 71974 82118 71986 82170
rect 72038 82118 72050 82170
rect 72102 82118 72114 82170
rect 72166 82118 74980 82170
rect 65320 82096 74980 82118
rect 63236 81784 63264 82052
rect 64874 81784 64880 81796
rect 63236 81756 64880 81784
rect 64874 81744 64880 81756
rect 64932 81744 64938 81796
rect 65320 81626 74980 81648
rect 65320 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74980 81626
rect 65320 81552 74980 81574
rect 65320 81082 74980 81104
rect 63236 80968 63264 81076
rect 65320 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 74980 81082
rect 65320 81008 74980 81030
rect 67082 80968 67088 80980
rect 63236 80940 67088 80968
rect 67082 80928 67088 80940
rect 67140 80928 67146 80980
rect 69750 80832 69756 80844
rect 63236 80804 69756 80832
rect 69750 80792 69756 80804
rect 69808 80792 69814 80844
rect 65320 80538 74980 80560
rect 65320 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74980 80538
rect 65320 80464 74980 80486
rect 65320 79994 74980 80016
rect 65320 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 74980 79994
rect 65320 79920 74980 79942
rect 64874 79880 64880 79892
rect 63236 79852 64880 79880
rect 64874 79840 64880 79852
rect 64932 79840 64938 79892
rect 65320 79450 74980 79472
rect 65320 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74980 79450
rect 65320 79376 74980 79398
rect 65320 78906 74980 78928
rect 63236 78724 63264 78896
rect 65320 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 74980 78906
rect 65320 78832 74980 78854
rect 66438 78724 66444 78736
rect 63236 78696 66444 78724
rect 66438 78684 66444 78696
rect 66496 78684 66502 78736
rect 69934 78656 69940 78668
rect 63236 78628 69940 78656
rect 69934 78616 69940 78628
rect 69992 78616 69998 78668
rect 65320 78362 74980 78384
rect 65320 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74980 78362
rect 65320 78288 74980 78310
rect 65320 77818 74980 77840
rect 65320 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 74980 77818
rect 65320 77744 74980 77766
rect 64874 77704 64880 77716
rect 63236 77676 64880 77704
rect 64874 77664 64880 77676
rect 64932 77664 64938 77716
rect 65320 77274 74980 77296
rect 65320 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74980 77274
rect 65320 77200 74980 77222
rect 65320 76730 74980 76752
rect 63236 76548 63264 76716
rect 65320 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 74980 76730
rect 65320 76656 74980 76678
rect 66254 76548 66260 76560
rect 63236 76520 66260 76548
rect 66254 76508 66260 76520
rect 66312 76508 66318 76560
rect 68462 76480 68468 76492
rect 63236 76452 68468 76480
rect 68462 76440 68468 76452
rect 68520 76440 68526 76492
rect 65320 76186 74980 76208
rect 65320 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74980 76186
rect 65320 76112 74980 76134
rect 65320 75642 74980 75664
rect 65320 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 74980 75642
rect 65320 75568 74980 75590
rect 63236 75188 63264 75512
rect 64874 75188 64880 75200
rect 63236 75160 64880 75188
rect 64874 75148 64880 75160
rect 64932 75148 64938 75200
rect 65320 75098 74980 75120
rect 65320 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74980 75098
rect 65320 75024 74980 75046
rect 67818 74644 67824 74656
rect 63236 74616 67824 74644
rect 63236 74536 63264 74616
rect 67818 74604 67824 74616
rect 67876 74604 67882 74656
rect 65320 74554 74980 74576
rect 65320 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 74980 74554
rect 65320 74480 74980 74502
rect 63236 74100 63264 74284
rect 66162 74100 66168 74112
rect 63236 74072 66168 74100
rect 66162 74060 66168 74072
rect 66220 74060 66226 74112
rect 65320 74010 74980 74032
rect 65320 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74980 74010
rect 65320 73936 74980 73958
rect 65320 73466 74980 73488
rect 65320 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 74980 73466
rect 65320 73392 74980 73414
rect 63236 73216 63264 73332
rect 64874 73216 64880 73228
rect 63236 73188 64880 73216
rect 64874 73176 64880 73188
rect 64932 73176 64938 73228
rect 65320 72922 74980 72944
rect 65320 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74980 72922
rect 65320 72848 74980 72870
rect 65320 72378 74980 72400
rect 63236 72196 63264 72356
rect 65320 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 74980 72378
rect 65320 72304 74980 72326
rect 66622 72196 66628 72208
rect 63236 72168 66628 72196
rect 66622 72156 66628 72168
rect 66680 72156 66686 72208
rect 63236 71788 63264 72104
rect 65320 71834 74980 71856
rect 65058 71788 65064 71800
rect 63236 71760 65064 71788
rect 65058 71748 65064 71760
rect 65116 71748 65122 71800
rect 65320 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74980 71834
rect 65320 71760 74980 71782
rect 65320 71290 74980 71312
rect 65320 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 74980 71290
rect 65320 71216 74980 71238
rect 63236 71148 63816 71176
rect 63788 71108 63816 71148
rect 64874 71108 64880 71120
rect 63788 71080 64880 71108
rect 64874 71068 64880 71080
rect 64932 71068 64938 71120
rect 65320 70746 74980 70768
rect 65320 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74980 70746
rect 65320 70672 74980 70694
rect 65320 70202 74980 70224
rect 63236 70020 63264 70176
rect 65320 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 74980 70202
rect 65320 70128 74980 70150
rect 65518 70020 65524 70032
rect 63236 69992 65524 70020
rect 65518 69980 65524 69992
rect 65576 69980 65582 70032
rect 63236 69612 63264 69924
rect 65320 69658 74980 69680
rect 63678 69612 63684 69624
rect 63236 69584 63684 69612
rect 63678 69572 63684 69584
rect 63736 69572 63742 69624
rect 65320 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74980 69658
rect 65320 69584 74980 69606
rect 65320 69114 74980 69136
rect 65320 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 74980 69114
rect 65320 69040 74980 69062
rect 63144 68972 63816 69000
rect 63788 68932 63816 68972
rect 64874 68932 64880 68944
rect 63788 68904 64880 68932
rect 64874 68892 64880 68904
rect 64932 68932 64938 68944
rect 66530 68932 66536 68944
rect 64932 68904 66536 68932
rect 64932 68892 64938 68904
rect 66530 68892 66536 68904
rect 66588 68892 66594 68944
rect 65320 68570 74980 68592
rect 65320 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74980 68570
rect 65320 68496 74980 68518
rect 65320 68026 74980 68048
rect 63236 67844 63264 67996
rect 65320 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 74980 68026
rect 65320 67952 74980 67974
rect 65886 67844 65892 67856
rect 63236 67816 65892 67844
rect 65886 67804 65892 67816
rect 65944 67804 65950 67856
rect 63494 67758 63500 67770
rect 63250 67730 63500 67758
rect 63494 67718 63500 67730
rect 63552 67718 63558 67770
rect 65320 67482 74980 67504
rect 65320 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74980 67482
rect 65320 67408 74980 67430
rect 65320 66938 74980 66960
rect 65320 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 74980 66938
rect 65320 66864 74980 66886
rect 63236 66484 63264 66792
rect 64874 66484 64880 66496
rect 63236 66456 64880 66484
rect 64874 66444 64880 66456
rect 64932 66444 64938 66496
rect 65320 66394 74980 66416
rect 65320 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74980 66394
rect 65320 66320 74980 66342
rect 65320 65850 74980 65872
rect 63236 65668 63264 65816
rect 65320 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 74980 65850
rect 65320 65776 74980 65798
rect 65426 65668 65432 65680
rect 63236 65640 65432 65668
rect 65426 65628 65432 65640
rect 65484 65628 65490 65680
rect 70394 65600 70400 65612
rect 63236 65572 70400 65600
rect 63236 65564 63264 65572
rect 70394 65560 70400 65572
rect 70452 65560 70458 65612
rect 65320 65306 74980 65328
rect 65320 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74980 65306
rect 65320 65232 74980 65254
rect 65320 64762 74980 64784
rect 65320 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 74980 64762
rect 65320 64688 74980 64710
rect 63236 64308 63264 64612
rect 64874 64308 64880 64320
rect 63236 64280 64880 64308
rect 64874 64268 64880 64280
rect 64932 64268 64938 64320
rect 65320 64218 74980 64240
rect 65320 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74980 64218
rect 65320 64144 74980 64166
rect 65320 63674 74980 63696
rect 63236 63560 63264 63636
rect 65320 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 74980 63674
rect 65320 63600 74980 63622
rect 65334 63560 65340 63572
rect 63236 63532 65340 63560
rect 65334 63520 65340 63532
rect 65392 63520 65398 63572
rect 63236 63220 63264 63384
rect 65702 63220 65708 63232
rect 63236 63192 65708 63220
rect 65702 63180 65708 63192
rect 65760 63180 65766 63232
rect 65320 63130 74980 63152
rect 65320 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74980 63130
rect 65320 63056 74980 63078
rect 65320 62586 74980 62608
rect 65320 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 74980 62586
rect 65320 62512 74980 62534
rect 63236 62132 63264 62432
rect 64874 62132 64880 62144
rect 63236 62104 64880 62132
rect 64874 62092 64880 62104
rect 64932 62092 64938 62144
rect 65320 62042 74980 62064
rect 65320 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74980 62042
rect 65320 61968 74980 61990
rect 65320 61498 74980 61520
rect 63236 61316 63264 61456
rect 65320 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 74980 61498
rect 65320 61424 74980 61446
rect 66070 61316 66076 61328
rect 63236 61288 66076 61316
rect 66070 61276 66076 61288
rect 66128 61276 66134 61328
rect 63236 60908 63264 61204
rect 65320 60954 74980 60976
rect 63586 60908 63592 60920
rect 63236 60880 63592 60908
rect 63586 60868 63592 60880
rect 63644 60868 63650 60920
rect 65320 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74980 60954
rect 65320 60880 74980 60902
rect 65320 60410 74980 60432
rect 65320 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 74980 60410
rect 65320 60336 74980 60358
rect 64874 60296 64880 60308
rect 63144 60268 64880 60296
rect 63144 60252 63172 60268
rect 64874 60256 64880 60268
rect 64932 60256 64938 60308
rect 65320 59866 74980 59888
rect 65320 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74980 59866
rect 65320 59792 74980 59814
rect 65320 59322 74980 59344
rect 63236 59140 63264 59276
rect 65320 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 74980 59322
rect 65320 59248 74980 59270
rect 65150 59140 65156 59152
rect 63236 59112 65156 59140
rect 65150 59100 65156 59112
rect 65208 59100 65214 59152
rect 69014 59072 69020 59084
rect 63236 59044 69020 59072
rect 63236 59024 63264 59044
rect 69014 59032 69020 59044
rect 69072 59032 69078 59084
rect 65320 58778 74980 58800
rect 65320 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74980 58778
rect 65320 58704 74980 58726
rect 65320 58234 74980 58256
rect 65320 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 74980 58234
rect 65320 58160 74980 58182
rect 63236 58052 63264 58072
rect 64874 58052 64880 58064
rect 63236 58024 64880 58052
rect 64874 58012 64880 58024
rect 64932 58012 64938 58064
rect 65320 57690 74980 57712
rect 65320 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74980 57690
rect 65320 57616 74980 57638
rect 65320 57146 74980 57168
rect 63236 56964 63264 57096
rect 65320 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 74980 57146
rect 65320 57072 74980 57094
rect 67542 56964 67548 56976
rect 63236 56936 67548 56964
rect 67542 56924 67548 56936
rect 67600 56924 67606 56976
rect 70486 56896 70492 56908
rect 63604 56868 70492 56896
rect 63604 56858 63632 56868
rect 63250 56830 63632 56858
rect 70486 56856 70492 56868
rect 70544 56856 70550 56908
rect 65320 56602 74980 56624
rect 65320 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74980 56602
rect 65320 56528 74980 56550
rect 65320 56058 74980 56080
rect 65320 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 74980 56058
rect 65320 55984 74980 56006
rect 63236 55604 63264 55892
rect 64874 55604 64880 55616
rect 63236 55576 64880 55604
rect 64874 55564 64880 55576
rect 64932 55564 64938 55616
rect 65320 55514 74980 55536
rect 65320 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74980 55514
rect 65320 55440 74980 55462
rect 65320 54970 74980 54992
rect 65320 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 74980 54970
rect 63236 54856 63264 54916
rect 65320 54896 74980 54918
rect 67726 54856 67732 54868
rect 63236 54828 67732 54856
rect 67726 54816 67732 54828
rect 67784 54816 67790 54868
rect 63236 54516 63264 54664
rect 65978 54516 65984 54528
rect 63236 54488 65984 54516
rect 65978 54476 65984 54488
rect 66036 54476 66042 54528
rect 65320 54426 74980 54448
rect 65320 54374 74210 54426
rect 74262 54374 74274 54426
rect 74326 54374 74338 54426
rect 74390 54374 74402 54426
rect 74454 54374 74466 54426
rect 74518 54374 74980 54426
rect 65320 54352 74980 54374
rect 65320 53882 74980 53904
rect 65320 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 74980 53882
rect 65320 53808 74980 53830
rect 63236 53564 63264 53712
rect 64874 53564 64880 53576
rect 63236 53536 64880 53564
rect 64874 53524 64880 53536
rect 64932 53524 64938 53576
rect 63236 53156 63264 53432
rect 65320 53338 74980 53360
rect 65320 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74980 53338
rect 65320 53264 74980 53286
rect 66898 53156 66904 53168
rect 63236 53128 66904 53156
rect 66898 53116 66904 53128
rect 66956 53116 66962 53168
rect 65320 52794 74980 52816
rect 65320 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 74980 52794
rect 63236 52612 63264 52736
rect 65320 52720 74980 52742
rect 66806 52612 66812 52624
rect 63236 52584 66812 52612
rect 66806 52572 66812 52584
rect 66864 52572 66870 52624
rect 63144 52476 63172 52484
rect 63770 52476 63776 52488
rect 63144 52448 63776 52476
rect 63770 52436 63776 52448
rect 63828 52436 63834 52488
rect 65610 52436 65616 52488
rect 65668 52436 65674 52488
rect 65889 52479 65947 52485
rect 65889 52445 65901 52479
rect 65935 52445 65947 52479
rect 65889 52439 65947 52445
rect 65904 52408 65932 52439
rect 63236 52380 65932 52408
rect 63236 52171 63264 52380
rect 65320 52250 74980 52272
rect 65320 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74980 52250
rect 65320 52176 74980 52198
rect 65610 52136 65616 52148
rect 63604 52108 65616 52136
rect 63250 52080 63632 52108
rect 65610 52096 65616 52108
rect 65668 52096 65674 52148
rect 65320 51706 74980 51728
rect 65320 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 74980 51706
rect 65320 51632 74980 51654
rect 63236 51524 63264 51532
rect 64874 51524 64880 51536
rect 63236 51496 64880 51524
rect 64874 51484 64880 51496
rect 64932 51524 64938 51536
rect 66346 51524 66352 51536
rect 64932 51496 66352 51524
rect 64932 51484 64938 51496
rect 66346 51484 66352 51496
rect 66404 51484 66410 51536
rect 65320 51162 74980 51184
rect 65320 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74980 51162
rect 65320 51088 74980 51110
rect 65320 50618 74980 50640
rect 65320 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 74980 50618
rect 63236 50504 63264 50556
rect 65320 50544 74980 50566
rect 67634 50504 67640 50516
rect 63236 50476 67640 50504
rect 67634 50464 67640 50476
rect 67692 50464 67698 50516
rect 63236 50300 63264 50304
rect 63770 50300 63776 50312
rect 63236 50272 63776 50300
rect 63770 50260 63776 50272
rect 63828 50260 63834 50312
rect 65613 50303 65671 50309
rect 65613 50300 65625 50303
rect 64846 50272 65625 50300
rect 64846 50232 64874 50272
rect 65613 50269 65625 50272
rect 65659 50269 65671 50303
rect 65613 50263 65671 50269
rect 63236 50204 64874 50232
rect 63236 49996 63264 50204
rect 65320 50074 74980 50096
rect 65320 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74980 50074
rect 65320 50000 74980 50022
rect 63250 49643 63632 49671
rect 63604 49620 63632 49643
rect 65613 49623 65671 49629
rect 65613 49620 65625 49623
rect 63604 49592 65625 49620
rect 65613 49589 65625 49592
rect 65659 49589 65671 49623
rect 65613 49583 65671 49589
rect 65320 49530 74980 49552
rect 65320 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 74980 49530
rect 65320 49456 74980 49478
rect 65613 49215 65671 49221
rect 65613 49181 65625 49215
rect 65659 49181 65671 49215
rect 65613 49175 65671 49181
rect 65242 49144 65248 49156
rect 63236 49116 65248 49144
rect 63236 48795 63264 49116
rect 65242 49104 65248 49116
rect 65300 49104 65306 49156
rect 65628 49076 65656 49175
rect 64846 49048 65656 49076
rect 64846 48736 64874 49048
rect 65320 48986 74980 49008
rect 65320 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74980 48986
rect 65320 48912 74980 48934
rect 63604 48729 64874 48736
rect 63250 48708 64874 48729
rect 63250 48701 63632 48708
rect 65320 48442 74980 48464
rect 65320 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 74980 48442
rect 65320 48368 74980 48390
rect 64966 48124 64972 48136
rect 63236 48096 64972 48124
rect 63236 48087 63264 48096
rect 64966 48084 64972 48096
rect 65024 48084 65030 48136
rect 63236 47716 63264 48007
rect 65320 47898 74980 47920
rect 65320 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74980 47898
rect 65320 47824 74980 47846
rect 64414 47716 64420 47728
rect 63236 47688 64420 47716
rect 64414 47676 64420 47688
rect 64472 47676 64478 47728
rect 63250 47376 63632 47393
rect 64598 47376 64604 47388
rect 63250 47365 64604 47376
rect 63604 47348 64604 47365
rect 64598 47336 64604 47348
rect 64656 47336 64662 47388
rect 65320 47354 74980 47376
rect 65320 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 74980 47354
rect 63236 47036 63264 47299
rect 65320 47280 74980 47302
rect 63862 47036 63868 47048
rect 63236 47008 63868 47036
rect 63862 46996 63868 47008
rect 63920 46996 63926 47048
rect 65613 47039 65671 47045
rect 65613 47005 65625 47039
rect 65659 47036 65671 47039
rect 68370 47036 68376 47048
rect 65659 47008 68376 47036
rect 65659 47005 65671 47008
rect 65613 46999 65671 47005
rect 68370 46996 68376 47008
rect 68428 46996 68434 47048
rect 65889 46971 65947 46977
rect 65889 46937 65901 46971
rect 65935 46968 65947 46971
rect 67174 46968 67180 46980
rect 65935 46940 67180 46968
rect 65935 46937 65947 46940
rect 65889 46931 65947 46937
rect 67174 46928 67180 46940
rect 67232 46928 67238 46980
rect 65320 46810 74980 46832
rect 65320 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74980 46810
rect 65320 46736 74980 46758
rect 65320 46266 74980 46288
rect 65320 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 74980 46266
rect 65320 46192 74980 46214
rect 63250 45949 63632 45977
rect 63604 45948 63632 45949
rect 64046 45948 64052 45960
rect 63604 45920 64052 45948
rect 64046 45908 64052 45920
rect 64104 45908 64110 45960
rect 63236 45744 63264 45883
rect 64138 45744 64144 45756
rect 63236 45716 64144 45744
rect 64138 45704 64144 45716
rect 64196 45704 64202 45756
rect 65320 45722 74980 45744
rect 65320 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74980 45722
rect 65320 45648 74980 45670
rect 63250 45268 63632 45269
rect 63954 45268 63960 45280
rect 63250 45241 63960 45268
rect 63604 45240 63960 45241
rect 63954 45228 63960 45240
rect 64012 45228 64018 45280
rect 65320 45178 74980 45200
rect 63236 44860 63264 45175
rect 65320 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 74980 45178
rect 65320 45104 74980 45126
rect 64966 44860 64972 44872
rect 63236 44832 64972 44860
rect 64966 44820 64972 44832
rect 65024 44820 65030 44872
rect 65320 44634 74980 44656
rect 65320 44582 74210 44634
rect 74262 44582 74274 44634
rect 74326 44582 74338 44634
rect 74390 44582 74402 44634
rect 74454 44582 74466 44634
rect 74518 44582 74980 44634
rect 63250 44533 63632 44561
rect 65320 44560 74980 44582
rect 63604 44520 63632 44533
rect 68186 44520 68192 44532
rect 63604 44492 68192 44520
rect 68186 44480 68192 44492
rect 68244 44480 68250 44532
rect 63236 44452 63264 44467
rect 68278 44452 68284 44464
rect 63236 44424 68284 44452
rect 68278 44412 68284 44424
rect 68336 44412 68342 44464
rect 65320 44090 74980 44112
rect 65320 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 74980 44090
rect 65320 44016 74980 44038
rect 64230 43840 64236 43852
rect 63236 43812 64236 43840
rect 64230 43800 64236 43812
rect 64288 43800 64294 43852
rect 65613 43775 65671 43781
rect 65613 43772 65625 43775
rect 63236 43744 65625 43772
rect 63236 43654 63264 43744
rect 65613 43741 65625 43744
rect 65659 43741 65671 43775
rect 65613 43735 65671 43741
rect 65320 43546 74980 43568
rect 65320 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74980 43546
rect 65320 43472 74980 43494
rect 63770 43296 63776 43308
rect 63236 43268 63776 43296
rect 63770 43256 63776 43268
rect 63828 43256 63834 43308
rect 68554 43092 68560 43104
rect 63512 43064 68560 43092
rect 63512 43032 63540 43064
rect 68554 43052 68560 43064
rect 68612 43052 68618 43104
rect 63250 43004 63540 43032
rect 65320 43002 74980 43024
rect 65320 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 74980 43002
rect 65320 42928 74980 42950
rect 66990 42712 66996 42764
rect 67048 42752 67054 42764
rect 68005 42755 68063 42761
rect 68005 42752 68017 42755
rect 67048 42724 68017 42752
rect 67048 42712 67054 42724
rect 68005 42721 68017 42724
rect 68051 42721 68063 42755
rect 68005 42715 68063 42721
rect 65613 42687 65671 42693
rect 65613 42684 65625 42687
rect 63236 42656 65625 42684
rect 63236 42402 63264 42656
rect 65613 42653 65625 42656
rect 65659 42653 65671 42687
rect 65613 42647 65671 42653
rect 68649 42687 68707 42693
rect 68649 42653 68661 42687
rect 68695 42684 68707 42687
rect 70026 42684 70032 42696
rect 68695 42656 70032 42684
rect 68695 42653 68707 42656
rect 68649 42647 68707 42653
rect 70026 42644 70032 42656
rect 70084 42644 70090 42696
rect 65320 42458 74980 42480
rect 65320 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74980 42458
rect 65320 42384 74980 42406
rect 63236 41732 63264 42042
rect 65320 41914 74980 41936
rect 65320 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 74980 41914
rect 65320 41840 74980 41862
rect 67082 41760 67088 41812
rect 67140 41760 67146 41812
rect 64874 41732 64880 41744
rect 63236 41704 64880 41732
rect 64874 41692 64880 41704
rect 64932 41692 64938 41744
rect 67729 41599 67787 41605
rect 67729 41565 67741 41599
rect 67775 41596 67787 41599
rect 70118 41596 70124 41608
rect 67775 41568 70124 41596
rect 67775 41565 67787 41568
rect 67729 41559 67787 41565
rect 70118 41556 70124 41568
rect 70176 41556 70182 41608
rect 65320 41370 74980 41392
rect 65320 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74980 41370
rect 65320 41296 74980 41318
rect 63236 40984 63264 41090
rect 65242 40984 65248 40996
rect 63236 40956 65248 40984
rect 65242 40944 65248 40956
rect 65300 40944 65306 40996
rect 68646 40916 68652 40928
rect 63512 40888 68652 40916
rect 63512 40852 63540 40888
rect 68646 40876 68652 40888
rect 68704 40876 68710 40928
rect 63250 40824 63540 40852
rect 65320 40826 74980 40848
rect 65320 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 74980 40826
rect 65320 40752 74980 40774
rect 66438 40672 66444 40724
rect 66496 40672 66502 40724
rect 67085 40511 67143 40517
rect 67085 40477 67097 40511
rect 67131 40508 67143 40511
rect 69198 40508 69204 40520
rect 67131 40480 69204 40508
rect 67131 40477 67143 40480
rect 67085 40471 67143 40477
rect 69198 40468 69204 40480
rect 69256 40468 69262 40520
rect 65320 40282 74980 40304
rect 65320 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74980 40282
rect 65320 40208 74980 40230
rect 63144 39868 63816 39896
rect 63144 39862 63172 39868
rect 63788 39828 63816 39868
rect 64874 39828 64880 39840
rect 63788 39800 64880 39828
rect 64874 39788 64880 39800
rect 64932 39788 64938 39840
rect 65320 39738 74980 39760
rect 65320 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 74980 39738
rect 65320 39664 74980 39686
rect 65613 39627 65671 39633
rect 65613 39593 65625 39627
rect 65659 39624 65671 39627
rect 66254 39624 66260 39636
rect 65659 39596 66260 39624
rect 65659 39593 65671 39596
rect 65613 39587 65671 39593
rect 66254 39584 66260 39596
rect 66312 39584 66318 39636
rect 66257 39423 66315 39429
rect 66257 39389 66269 39423
rect 66303 39420 66315 39423
rect 67450 39420 67456 39432
rect 66303 39392 67456 39420
rect 66303 39389 66315 39392
rect 66257 39383 66315 39389
rect 67450 39380 67456 39392
rect 67508 39380 67514 39432
rect 65320 39194 74980 39216
rect 65320 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74980 39194
rect 65320 39120 74980 39142
rect 63236 38808 63264 38910
rect 65242 38808 65248 38820
rect 63236 38780 65248 38808
rect 65242 38768 65248 38780
rect 65300 38768 65306 38820
rect 67910 38740 67916 38752
rect 63236 38712 67916 38740
rect 63236 38658 63264 38712
rect 67910 38700 67916 38712
rect 67968 38700 67974 38752
rect 65320 38650 74980 38672
rect 65320 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 74980 38650
rect 65320 38576 74980 38598
rect 65613 38539 65671 38545
rect 65613 38505 65625 38539
rect 65659 38536 65671 38539
rect 67818 38536 67824 38548
rect 65659 38508 67824 38536
rect 65659 38505 65671 38508
rect 65613 38499 65671 38505
rect 67818 38496 67824 38508
rect 67876 38496 67882 38548
rect 66257 38335 66315 38341
rect 66257 38301 66269 38335
rect 66303 38332 66315 38335
rect 66990 38332 66996 38344
rect 66303 38304 66996 38332
rect 66303 38301 66315 38304
rect 66257 38295 66315 38301
rect 66990 38292 66996 38304
rect 67048 38292 67054 38344
rect 65320 38106 74980 38128
rect 65320 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74980 38106
rect 65320 38032 74980 38054
rect 63236 37380 63264 37682
rect 65320 37562 74980 37584
rect 65320 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 74980 37562
rect 65320 37488 74980 37510
rect 64874 37380 64880 37392
rect 63236 37352 64880 37380
rect 64874 37340 64880 37352
rect 64932 37340 64938 37392
rect 66257 37247 66315 37253
rect 66257 37213 66269 37247
rect 66303 37244 66315 37247
rect 67266 37244 67272 37256
rect 66303 37216 67272 37244
rect 66303 37213 66315 37216
rect 66257 37207 66315 37213
rect 67266 37204 67272 37216
rect 67324 37204 67330 37256
rect 65613 37179 65671 37185
rect 65613 37145 65625 37179
rect 65659 37176 65671 37179
rect 66622 37176 66628 37188
rect 65659 37148 66628 37176
rect 65659 37145 65671 37148
rect 65613 37139 65671 37145
rect 66622 37136 66628 37148
rect 66680 37136 66686 37188
rect 65320 37018 74980 37040
rect 65320 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74980 37018
rect 65320 36944 74980 36966
rect 63236 36564 63264 36730
rect 65794 36564 65800 36576
rect 63236 36536 65800 36564
rect 65794 36524 65800 36536
rect 65852 36524 65858 36576
rect 63236 36360 63264 36478
rect 65320 36474 74980 36496
rect 65320 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 74980 36474
rect 65320 36400 74980 36422
rect 63236 36332 64874 36360
rect 64846 36292 64874 36332
rect 65518 36320 65524 36372
rect 65576 36360 65582 36372
rect 65613 36363 65671 36369
rect 65613 36360 65625 36363
rect 65576 36332 65625 36360
rect 65576 36320 65582 36332
rect 65613 36329 65625 36332
rect 65659 36329 65671 36363
rect 65613 36323 65671 36329
rect 68094 36292 68100 36304
rect 64846 36264 68100 36292
rect 68094 36252 68100 36264
rect 68152 36252 68158 36304
rect 66257 36159 66315 36165
rect 66257 36125 66269 36159
rect 66303 36156 66315 36159
rect 67358 36156 67364 36168
rect 66303 36128 67364 36156
rect 66303 36125 66315 36128
rect 66257 36119 66315 36125
rect 67358 36116 67364 36128
rect 67416 36116 67422 36168
rect 65320 35930 74980 35952
rect 65320 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74980 35930
rect 65320 35856 74980 35878
rect 66530 35708 66536 35760
rect 66588 35708 66594 35760
rect 65797 35683 65855 35689
rect 65797 35649 65809 35683
rect 65843 35680 65855 35683
rect 68002 35680 68008 35692
rect 65843 35652 68008 35680
rect 65843 35649 65855 35652
rect 65797 35643 65855 35649
rect 68002 35640 68008 35652
rect 68060 35640 68066 35692
rect 63236 35204 63264 35502
rect 65320 35386 74980 35408
rect 65320 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 74980 35386
rect 65320 35312 74980 35334
rect 65613 35275 65671 35281
rect 65613 35241 65625 35275
rect 65659 35272 65671 35275
rect 65886 35272 65892 35284
rect 65659 35244 65892 35272
rect 65659 35241 65671 35244
rect 65613 35235 65671 35241
rect 65886 35232 65892 35244
rect 65944 35232 65950 35284
rect 64874 35204 64880 35216
rect 63236 35176 64880 35204
rect 64874 35164 64880 35176
rect 64932 35164 64938 35216
rect 66257 35071 66315 35077
rect 66257 35037 66269 35071
rect 66303 35068 66315 35071
rect 66622 35068 66628 35080
rect 66303 35040 66628 35068
rect 66303 35037 66315 35040
rect 66257 35031 66315 35037
rect 66622 35028 66628 35040
rect 66680 35028 66686 35080
rect 65320 34842 74980 34864
rect 65320 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74980 34842
rect 65320 34768 74980 34790
rect 63250 34536 63632 34564
rect 63604 34524 63632 34536
rect 65242 34524 65248 34536
rect 63604 34496 65248 34524
rect 65242 34484 65248 34496
rect 65300 34484 65306 34536
rect 65320 34298 74980 34320
rect 63236 33980 63264 34298
rect 65320 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 74980 34298
rect 65320 34224 74980 34246
rect 66898 34144 66904 34196
rect 66956 34144 66962 34196
rect 64782 33980 64788 33992
rect 63236 33952 64788 33980
rect 64782 33940 64788 33952
rect 64840 33940 64846 33992
rect 65610 33872 65616 33924
rect 65668 33872 65674 33924
rect 65320 33754 74980 33776
rect 65320 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74980 33754
rect 65320 33680 74980 33702
rect 65426 33600 65432 33652
rect 65484 33640 65490 33652
rect 65613 33643 65671 33649
rect 65613 33640 65625 33643
rect 65484 33612 65625 33640
rect 65484 33600 65490 33612
rect 65613 33609 65625 33612
rect 65659 33609 65671 33643
rect 65613 33603 65671 33609
rect 66257 33439 66315 33445
rect 66257 33405 66269 33439
rect 66303 33436 66315 33439
rect 66714 33436 66720 33448
rect 66303 33408 66720 33436
rect 66303 33405 66315 33408
rect 66257 33399 66315 33405
rect 66714 33396 66720 33408
rect 66772 33396 66778 33448
rect 63236 33300 63264 33322
rect 64874 33300 64880 33312
rect 63236 33272 64880 33300
rect 64874 33260 64880 33272
rect 64932 33260 64938 33312
rect 65320 33210 74980 33232
rect 65320 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 74980 33210
rect 65320 33136 74980 33158
rect 65334 33056 65340 33108
rect 65392 33096 65398 33108
rect 65613 33099 65671 33105
rect 65613 33096 65625 33099
rect 65392 33068 65625 33096
rect 65392 33056 65398 33068
rect 65613 33065 65625 33068
rect 65659 33065 65671 33099
rect 65613 33059 65671 33065
rect 66438 32988 66444 33040
rect 66496 33028 66502 33040
rect 67542 33028 67548 33040
rect 66496 33000 67548 33028
rect 66496 32988 66502 33000
rect 67542 32988 67548 33000
rect 67600 32988 67606 33040
rect 66257 32895 66315 32901
rect 66257 32861 66269 32895
rect 66303 32892 66315 32895
rect 67542 32892 67548 32904
rect 66303 32864 67548 32892
rect 66303 32861 66315 32864
rect 66257 32855 66315 32861
rect 67542 32852 67548 32864
rect 67600 32852 67606 32904
rect 65320 32666 74980 32688
rect 65320 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74980 32666
rect 65320 32592 74980 32614
rect 63236 32212 63264 32370
rect 65334 32212 65340 32224
rect 63236 32184 65340 32212
rect 65334 32172 65340 32184
rect 65392 32172 65398 32224
rect 65320 32122 74980 32144
rect 63236 31804 63264 32118
rect 65320 32070 71858 32122
rect 71910 32070 71922 32122
rect 71974 32070 71986 32122
rect 72038 32070 72050 32122
rect 72102 32070 72114 32122
rect 72166 32070 74980 32122
rect 65320 32048 74980 32070
rect 65613 32011 65671 32017
rect 65613 31977 65625 32011
rect 65659 32008 65671 32011
rect 66070 32008 66076 32020
rect 65659 31980 66076 32008
rect 65659 31977 65671 31980
rect 65613 31971 65671 31977
rect 66070 31968 66076 31980
rect 66128 31968 66134 32020
rect 64414 31804 64420 31816
rect 63236 31776 64420 31804
rect 64414 31764 64420 31776
rect 64472 31764 64478 31816
rect 66257 31807 66315 31813
rect 66257 31773 66269 31807
rect 66303 31804 66315 31807
rect 67082 31804 67088 31816
rect 66303 31776 67088 31804
rect 66303 31773 66315 31776
rect 66257 31767 66315 31773
rect 67082 31764 67088 31776
rect 67140 31764 67146 31816
rect 65320 31578 74980 31600
rect 65320 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74980 31578
rect 65320 31504 74980 31526
rect 63236 31124 63264 31142
rect 64874 31124 64880 31136
rect 63236 31096 64880 31124
rect 64874 31084 64880 31096
rect 64932 31084 64938 31136
rect 65320 31034 74980 31056
rect 65320 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 74980 31034
rect 65320 30960 74980 30982
rect 65150 30880 65156 30932
rect 65208 30920 65214 30932
rect 65613 30923 65671 30929
rect 65613 30920 65625 30923
rect 65208 30892 65625 30920
rect 65208 30880 65214 30892
rect 65613 30889 65625 30892
rect 65659 30889 65671 30923
rect 65613 30883 65671 30889
rect 66257 30719 66315 30725
rect 66257 30685 66269 30719
rect 66303 30716 66315 30719
rect 66806 30716 66812 30728
rect 66303 30688 66812 30716
rect 66303 30685 66315 30688
rect 66257 30679 66315 30685
rect 66806 30676 66812 30688
rect 66864 30676 66870 30728
rect 65320 30490 74980 30512
rect 65320 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74980 30490
rect 65320 30416 74980 30438
rect 63236 30036 63264 30190
rect 65426 30036 65432 30048
rect 63236 30008 65432 30036
rect 65426 29996 65432 30008
rect 65484 29996 65490 30048
rect 65320 29946 74980 29968
rect 63236 29628 63264 29938
rect 65320 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 74980 29946
rect 65320 29872 74980 29894
rect 65613 29835 65671 29841
rect 65613 29801 65625 29835
rect 65659 29832 65671 29835
rect 66438 29832 66444 29844
rect 65659 29804 66444 29832
rect 65659 29801 65671 29804
rect 65613 29795 65671 29801
rect 66438 29792 66444 29804
rect 66496 29792 66502 29844
rect 64322 29628 64328 29640
rect 63236 29600 64328 29628
rect 64322 29588 64328 29600
rect 64380 29588 64386 29640
rect 66257 29631 66315 29637
rect 66257 29597 66269 29631
rect 66303 29628 66315 29631
rect 66438 29628 66444 29640
rect 66303 29600 66444 29628
rect 66303 29597 66315 29600
rect 66257 29591 66315 29597
rect 66438 29588 66444 29600
rect 66496 29588 66502 29640
rect 65320 29402 74980 29424
rect 65320 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74980 29402
rect 65320 29328 74980 29350
rect 63236 28676 63264 28962
rect 65320 28858 74980 28880
rect 65320 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 74980 28858
rect 65320 28784 74980 28806
rect 65613 28747 65671 28753
rect 65613 28713 65625 28747
rect 65659 28744 65671 28747
rect 67726 28744 67732 28756
rect 65659 28716 67732 28744
rect 65659 28713 65671 28716
rect 65613 28707 65671 28713
rect 67726 28704 67732 28716
rect 67784 28704 67790 28756
rect 64874 28676 64880 28688
rect 63236 28648 64880 28676
rect 64874 28636 64880 28648
rect 64932 28636 64938 28688
rect 66254 28500 66260 28552
rect 66312 28500 66318 28552
rect 65320 28314 74980 28336
rect 65320 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74980 28314
rect 65320 28240 74980 28262
rect 63236 27860 63264 28010
rect 65886 27860 65892 27872
rect 63236 27832 65892 27860
rect 65886 27820 65892 27832
rect 65944 27820 65950 27872
rect 65320 27770 74980 27792
rect 63236 27656 63264 27758
rect 65320 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 74980 27770
rect 65320 27696 74980 27718
rect 64506 27656 64512 27668
rect 63236 27628 64512 27656
rect 64506 27616 64512 27628
rect 64564 27616 64570 27668
rect 65613 27591 65671 27597
rect 65613 27557 65625 27591
rect 65659 27588 65671 27591
rect 66530 27588 66536 27600
rect 65659 27560 66536 27588
rect 65659 27557 65671 27560
rect 65613 27551 65671 27557
rect 66530 27548 66536 27560
rect 66588 27548 66594 27600
rect 66257 27455 66315 27461
rect 66257 27421 66269 27455
rect 66303 27452 66315 27455
rect 66990 27452 66996 27464
rect 66303 27424 66996 27452
rect 66303 27421 66315 27424
rect 66257 27415 66315 27421
rect 66990 27412 66996 27424
rect 67048 27412 67054 27464
rect 65320 27226 74980 27248
rect 65320 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74980 27226
rect 65320 27152 74980 27174
rect 64874 27044 64880 27056
rect 63236 27016 64880 27044
rect 63236 26782 63264 27016
rect 64874 27004 64880 27016
rect 64932 27044 64938 27056
rect 68830 27044 68836 27056
rect 64932 27016 68836 27044
rect 64932 27004 64938 27016
rect 68830 27004 68836 27016
rect 68888 27004 68894 27056
rect 65797 26979 65855 26985
rect 65797 26945 65809 26979
rect 65843 26976 65855 26979
rect 68738 26976 68744 26988
rect 65843 26948 68744 26976
rect 65843 26945 65855 26948
rect 65797 26939 65855 26945
rect 68738 26936 68744 26948
rect 68796 26936 68802 26988
rect 66346 26868 66352 26920
rect 66404 26868 66410 26920
rect 65320 26682 74980 26704
rect 65320 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 74980 26682
rect 65320 26608 74980 26630
rect 65613 26571 65671 26577
rect 65613 26537 65625 26571
rect 65659 26568 65671 26571
rect 67634 26568 67640 26580
rect 65659 26540 67640 26568
rect 65659 26537 65671 26540
rect 65613 26531 65671 26537
rect 67634 26528 67640 26540
rect 67692 26528 67698 26580
rect 66257 26367 66315 26373
rect 66257 26333 66269 26367
rect 66303 26364 66315 26367
rect 66530 26364 66536 26376
rect 66303 26336 66536 26364
rect 66303 26333 66315 26336
rect 66257 26327 66315 26333
rect 66530 26324 66536 26336
rect 66588 26324 66594 26376
rect 65320 26138 74980 26160
rect 65320 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74980 26138
rect 65320 26064 74980 26086
rect 63236 25684 63264 25830
rect 65610 25684 65616 25696
rect 63236 25656 65616 25684
rect 65610 25644 65616 25656
rect 65668 25644 65674 25696
rect 65320 25594 74980 25616
rect 63236 25276 63264 25578
rect 65320 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 74980 25594
rect 65320 25520 74980 25542
rect 63770 25276 63776 25288
rect 63236 25248 63776 25276
rect 63770 25236 63776 25248
rect 63828 25236 63834 25288
rect 65320 25050 74980 25072
rect 65320 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74980 25050
rect 65320 24976 74980 24998
rect 63236 24324 63264 24602
rect 65320 24506 74980 24528
rect 65320 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 74980 24506
rect 65320 24432 74980 24454
rect 65613 24395 65671 24401
rect 65613 24361 65625 24395
rect 65659 24392 65671 24395
rect 68278 24392 68284 24404
rect 65659 24364 68284 24392
rect 65659 24361 65671 24364
rect 65613 24355 65671 24361
rect 68278 24352 68284 24364
rect 68336 24352 68342 24404
rect 65150 24324 65156 24336
rect 63236 24296 65156 24324
rect 65150 24284 65156 24296
rect 65208 24284 65214 24336
rect 66257 24191 66315 24197
rect 66257 24157 66269 24191
rect 66303 24188 66315 24191
rect 66346 24188 66352 24200
rect 66303 24160 66352 24188
rect 66303 24157 66315 24160
rect 66257 24151 66315 24157
rect 66346 24148 66352 24160
rect 66404 24148 66410 24200
rect 65320 23962 74980 23984
rect 65320 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74980 23962
rect 65320 23888 74980 23910
rect 64966 23808 64972 23860
rect 65024 23848 65030 23860
rect 65613 23851 65671 23857
rect 65613 23848 65625 23851
rect 65024 23820 65625 23848
rect 65024 23808 65030 23820
rect 65613 23817 65625 23820
rect 65659 23817 65671 23851
rect 65613 23811 65671 23817
rect 66530 23740 66536 23792
rect 66588 23780 66594 23792
rect 66990 23780 66996 23792
rect 66588 23752 66996 23780
rect 66588 23740 66594 23752
rect 66990 23740 66996 23752
rect 67048 23740 67054 23792
rect 63236 23508 63264 23650
rect 66257 23647 66315 23653
rect 66257 23613 66269 23647
rect 66303 23644 66315 23647
rect 66530 23644 66536 23656
rect 66303 23616 66536 23644
rect 66303 23613 66315 23616
rect 66257 23607 66315 23613
rect 66530 23604 66536 23616
rect 66588 23604 66594 23656
rect 66070 23508 66076 23520
rect 63236 23480 66076 23508
rect 66070 23468 66076 23480
rect 66128 23468 66134 23520
rect 65320 23418 74980 23440
rect 63236 23304 63264 23398
rect 65320 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 74980 23418
rect 65320 23344 74980 23366
rect 65613 23307 65671 23313
rect 63236 23276 64874 23304
rect 64846 23236 64874 23276
rect 65613 23273 65625 23307
rect 65659 23304 65671 23307
rect 68186 23304 68192 23316
rect 65659 23276 68192 23304
rect 65659 23273 65671 23276
rect 65613 23267 65671 23273
rect 68186 23264 68192 23276
rect 68244 23264 68250 23316
rect 68922 23236 68928 23248
rect 64846 23208 68928 23236
rect 68922 23196 68928 23208
rect 68980 23196 68986 23248
rect 66257 23103 66315 23109
rect 66257 23069 66269 23103
rect 66303 23100 66315 23103
rect 66530 23100 66536 23112
rect 66303 23072 66536 23100
rect 66303 23069 66315 23072
rect 66257 23063 66315 23069
rect 66530 23060 66536 23072
rect 66588 23060 66594 23112
rect 65320 22874 74980 22896
rect 65320 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74980 22874
rect 65320 22800 74980 22822
rect 63236 22148 63264 22422
rect 65320 22330 74980 22352
rect 65320 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 74980 22330
rect 65320 22256 74980 22278
rect 65150 22148 65156 22160
rect 63236 22120 65156 22148
rect 65150 22108 65156 22120
rect 65208 22108 65214 22160
rect 65320 21786 74980 21808
rect 65320 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74980 21786
rect 65320 21712 74980 21734
rect 70578 21536 70584 21548
rect 63604 21508 70584 21536
rect 63604 21484 63632 21508
rect 70578 21496 70584 21508
rect 70636 21496 70642 21548
rect 63250 21456 63632 21484
rect 65320 21242 74980 21264
rect 63236 21128 63264 21218
rect 65320 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 74980 21242
rect 65320 21168 74980 21190
rect 67818 21128 67824 21140
rect 63236 21100 67824 21128
rect 67818 21088 67824 21100
rect 67876 21088 67882 21140
rect 65320 20698 74980 20720
rect 65320 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74980 20698
rect 65320 20624 74980 20646
rect 65150 20244 65156 20256
rect 63236 20216 65156 20244
rect 65150 20204 65156 20216
rect 65208 20204 65214 20256
rect 65320 20154 74980 20176
rect 65320 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 74980 20154
rect 65320 20080 74980 20102
rect 65320 19610 74980 19632
rect 65320 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74980 19610
rect 65320 19536 74980 19558
rect 63236 19156 63264 19290
rect 65518 19156 65524 19168
rect 63236 19128 65524 19156
rect 65518 19116 65524 19128
rect 65576 19116 65582 19168
rect 65320 19066 74980 19088
rect 63236 18748 63264 19038
rect 65320 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 74980 19066
rect 65320 18992 74980 19014
rect 64690 18748 64696 18760
rect 63236 18720 64696 18748
rect 64690 18708 64696 18720
rect 64748 18708 64754 18760
rect 65320 18522 74980 18544
rect 65320 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74980 18522
rect 65320 18448 74980 18470
rect 63236 18000 63264 18062
rect 65150 18000 65156 18012
rect 63236 17972 65156 18000
rect 65150 17960 65156 17972
rect 65208 17960 65214 18012
rect 65320 17978 74980 18000
rect 65320 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 74980 17978
rect 65320 17904 74980 17926
rect 65320 17434 74980 17456
rect 65320 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74980 17434
rect 65320 17360 74980 17382
rect 70670 17184 70676 17196
rect 63604 17156 70676 17184
rect 63604 17124 63632 17156
rect 70670 17144 70676 17156
rect 70728 17144 70734 17196
rect 63250 17096 63632 17124
rect 65320 16890 74980 16912
rect 63236 16640 63264 16858
rect 65320 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 74980 16890
rect 65320 16816 74980 16838
rect 63236 16612 63724 16640
rect 63696 16584 63724 16612
rect 63678 16532 63684 16584
rect 63736 16532 63742 16584
rect 65320 16346 74980 16368
rect 65320 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74980 16346
rect 65320 16272 74980 16294
rect 63236 15620 63264 15882
rect 65320 15802 74980 15824
rect 65320 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 74980 15802
rect 65320 15728 74980 15750
rect 65150 15620 65156 15632
rect 63236 15592 65156 15620
rect 65150 15580 65156 15592
rect 65208 15580 65214 15632
rect 65320 15258 74980 15280
rect 65320 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74980 15258
rect 65320 15184 74980 15206
rect 63236 14804 63264 14930
rect 65518 14804 65524 14816
rect 63236 14776 65524 14804
rect 65518 14764 65524 14776
rect 65576 14764 65582 14816
rect 65320 14714 74980 14736
rect 63236 14600 63264 14678
rect 65320 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 74980 14714
rect 65320 14640 74980 14662
rect 67634 14600 67640 14612
rect 63236 14572 67640 14600
rect 67634 14560 67640 14572
rect 67692 14560 67698 14612
rect 65320 14170 74980 14192
rect 65320 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74980 14170
rect 65320 14096 74980 14118
rect 65150 13716 65156 13728
rect 63250 13688 65156 13716
rect 65150 13676 65156 13688
rect 65208 13676 65214 13728
rect 65320 13626 74980 13648
rect 65320 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 74980 13626
rect 65320 13552 74980 13574
rect 65320 13082 74980 13104
rect 65320 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74980 13082
rect 65320 13008 74980 13030
rect 64874 12764 64880 12776
rect 63250 12736 64880 12764
rect 64874 12724 64880 12736
rect 64932 12724 64938 12776
rect 67726 12628 67732 12640
rect 63236 12600 67732 12628
rect 63236 12498 63264 12600
rect 67726 12588 67732 12600
rect 67784 12588 67790 12640
rect 65320 12538 74980 12560
rect 65320 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 74980 12538
rect 65320 12464 74980 12486
rect 63954 12248 63960 12300
rect 64012 12288 64018 12300
rect 64690 12288 64696 12300
rect 64012 12260 64696 12288
rect 64012 12248 64018 12260
rect 64690 12248 64696 12260
rect 64748 12248 64754 12300
rect 65320 11994 74980 12016
rect 65320 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74980 11994
rect 65320 11920 74980 11942
rect 63236 11268 63264 11522
rect 65320 11450 74980 11472
rect 65320 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 74980 11450
rect 65320 11376 74980 11398
rect 64598 11296 64604 11348
rect 64656 11336 64662 11348
rect 64782 11336 64788 11348
rect 64656 11308 64788 11336
rect 64656 11296 64662 11308
rect 64782 11296 64788 11308
rect 64840 11296 64846 11348
rect 65150 11268 65156 11280
rect 63236 11240 65156 11268
rect 65150 11228 65156 11240
rect 65208 11268 65214 11280
rect 65334 11268 65340 11280
rect 65208 11240 65340 11268
rect 65208 11228 65214 11240
rect 65334 11228 65340 11240
rect 65392 11228 65398 11280
rect 64230 11160 64236 11212
rect 64288 11200 64294 11212
rect 64598 11200 64604 11212
rect 64288 11172 64604 11200
rect 64288 11160 64294 11172
rect 64598 11160 64604 11172
rect 64656 11160 64662 11212
rect 64230 11024 64236 11076
rect 64288 11064 64294 11076
rect 67174 11064 67180 11076
rect 64288 11036 67180 11064
rect 64288 11024 64294 11036
rect 67174 11024 67180 11036
rect 67232 11024 67238 11076
rect 65320 10906 74980 10928
rect 65320 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74980 10906
rect 65320 10832 74980 10854
rect 63236 10452 63264 10570
rect 64874 10548 64880 10600
rect 64932 10588 64938 10600
rect 65150 10588 65156 10600
rect 64932 10560 65156 10588
rect 64932 10548 64938 10560
rect 65150 10548 65156 10560
rect 65208 10548 65214 10600
rect 64874 10452 64880 10464
rect 63236 10424 64880 10452
rect 64874 10412 64880 10424
rect 64932 10412 64938 10464
rect 65320 10362 74980 10384
rect 63402 10332 63408 10344
rect 63250 10304 63408 10332
rect 63402 10292 63408 10304
rect 63460 10292 63466 10344
rect 65320 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 74980 10362
rect 65320 10288 74980 10310
rect 65320 9818 74980 9840
rect 65320 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74980 9818
rect 65320 9744 74980 9766
rect 63236 9160 63264 9342
rect 65320 9274 74980 9296
rect 65320 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 74980 9274
rect 65320 9200 74980 9222
rect 65334 9160 65340 9172
rect 63236 9132 65340 9160
rect 65334 9120 65340 9132
rect 65392 9120 65398 9172
rect 65320 8730 74980 8752
rect 65320 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74980 8730
rect 65320 8656 74980 8678
rect 65320 8186 74980 8208
rect 65320 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 74980 8186
rect 65320 8112 74980 8134
rect 64230 7936 64236 7948
rect 60706 7908 64236 7936
rect 59554 7760 59560 7812
rect 59612 7800 59618 7812
rect 60706 7800 60734 7908
rect 64230 7896 64236 7908
rect 64288 7896 64294 7948
rect 61654 7828 61660 7880
rect 61712 7868 61718 7880
rect 63494 7868 63500 7880
rect 61712 7840 63500 7868
rect 61712 7828 61718 7840
rect 63494 7828 63500 7840
rect 63552 7828 63558 7880
rect 59612 7772 60734 7800
rect 59612 7760 59618 7772
rect 62482 7760 62488 7812
rect 62540 7800 62546 7812
rect 64966 7800 64972 7812
rect 62540 7772 64972 7800
rect 62540 7760 62546 7772
rect 64966 7760 64972 7772
rect 65024 7760 65030 7812
rect 52270 7692 52276 7744
rect 52328 7732 52334 7744
rect 63678 7732 63684 7744
rect 52328 7704 63684 7732
rect 52328 7692 52334 7704
rect 63678 7692 63684 7704
rect 63736 7692 63742 7744
rect 56134 7624 56140 7676
rect 56192 7664 56198 7676
rect 63402 7664 63408 7676
rect 56192 7636 63408 7664
rect 56192 7624 56198 7636
rect 63402 7624 63408 7636
rect 63460 7624 63466 7676
rect 65320 7642 74980 7664
rect 56502 7556 56508 7608
rect 56560 7596 56566 7608
rect 63586 7596 63592 7608
rect 56560 7568 63592 7596
rect 56560 7556 56566 7568
rect 63586 7556 63592 7568
rect 63644 7556 63650 7608
rect 65320 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74980 7642
rect 65320 7568 74980 7590
rect 48222 7488 48228 7540
rect 48280 7528 48286 7540
rect 64322 7528 64328 7540
rect 48280 7500 64328 7528
rect 48280 7488 48286 7500
rect 64322 7488 64328 7500
rect 64380 7488 64386 7540
rect 59170 7420 59176 7472
rect 59228 7460 59234 7472
rect 68370 7460 68376 7472
rect 59228 7432 68376 7460
rect 59228 7420 59234 7432
rect 68370 7420 68376 7432
rect 68428 7420 68434 7472
rect 62758 7352 62764 7404
rect 62816 7392 62822 7404
rect 65702 7392 65708 7404
rect 62816 7364 65708 7392
rect 62816 7352 62822 7364
rect 65702 7352 65708 7364
rect 65760 7352 65766 7404
rect 63034 7284 63040 7336
rect 63092 7324 63098 7336
rect 65518 7324 65524 7336
rect 63092 7296 65524 7324
rect 63092 7284 63098 7296
rect 65518 7284 65524 7296
rect 65576 7284 65582 7336
rect 60366 7216 60372 7268
rect 60424 7256 60430 7268
rect 64690 7256 64696 7268
rect 60424 7228 64696 7256
rect 60424 7216 60430 7228
rect 64690 7216 64696 7228
rect 64748 7216 64754 7268
rect 65320 7098 74980 7120
rect 60090 7012 60096 7064
rect 60148 7052 60154 7064
rect 65150 7052 65156 7064
rect 60148 7024 65156 7052
rect 60148 7012 60154 7024
rect 65150 7012 65156 7024
rect 65208 7012 65214 7064
rect 65320 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 74980 7098
rect 65320 7024 74980 7046
rect 55582 6944 55588 6996
rect 55640 6984 55646 6996
rect 55640 6956 60136 6984
rect 55640 6944 55646 6956
rect 55674 6876 55680 6928
rect 55732 6916 55738 6928
rect 55732 6888 56180 6916
rect 55732 6876 55738 6888
rect 48866 6808 48872 6860
rect 48924 6848 48930 6860
rect 56042 6848 56048 6860
rect 48924 6820 56048 6848
rect 48924 6808 48930 6820
rect 56042 6808 56048 6820
rect 56100 6808 56106 6860
rect 56152 6848 56180 6888
rect 59998 6848 60004 6860
rect 56152 6820 60004 6848
rect 59998 6808 60004 6820
rect 60056 6808 60062 6860
rect 60108 6848 60136 6956
rect 65720 6888 66760 6916
rect 65720 6848 65748 6888
rect 60108 6820 65748 6848
rect 65794 6808 65800 6860
rect 65852 6848 65858 6860
rect 66622 6848 66628 6860
rect 65852 6820 66628 6848
rect 65852 6808 65858 6820
rect 66622 6808 66628 6820
rect 66680 6808 66686 6860
rect 66732 6848 66760 6888
rect 68922 6848 68928 6860
rect 66732 6820 68928 6848
rect 68922 6808 68928 6820
rect 68980 6808 68986 6860
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 64874 6780 64880 6792
rect 27580 6752 64880 6780
rect 27580 6740 27586 6752
rect 64874 6740 64880 6752
rect 64932 6740 64938 6792
rect 65150 6740 65156 6792
rect 65208 6780 65214 6792
rect 66806 6780 66812 6792
rect 65208 6752 66812 6780
rect 65208 6740 65214 6752
rect 66806 6740 66812 6752
rect 66864 6740 66870 6792
rect 23290 6672 23296 6724
rect 23348 6712 23354 6724
rect 70670 6712 70676 6724
rect 23348 6684 70676 6712
rect 23348 6672 23354 6684
rect 70670 6672 70676 6684
rect 70728 6672 70734 6724
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 70578 6644 70584 6656
rect 24820 6616 70584 6644
rect 24820 6604 24826 6616
rect 70578 6604 70584 6616
rect 70636 6604 70642 6656
rect 25866 6536 25872 6588
rect 25924 6576 25930 6588
rect 62482 6576 62488 6588
rect 25924 6548 62488 6576
rect 25924 6536 25930 6548
rect 62482 6536 62488 6548
rect 62540 6536 62546 6588
rect 63494 6536 63500 6588
rect 63552 6576 63558 6588
rect 64966 6576 64972 6588
rect 63552 6548 64972 6576
rect 63552 6536 63558 6548
rect 64966 6536 64972 6548
rect 65024 6536 65030 6588
rect 65320 6554 74980 6576
rect 28626 6468 28632 6520
rect 28684 6508 28690 6520
rect 46382 6508 46388 6520
rect 28684 6480 46388 6508
rect 28684 6468 28690 6480
rect 46382 6468 46388 6480
rect 46440 6468 46446 6520
rect 54662 6468 54668 6520
rect 54720 6508 54726 6520
rect 59538 6508 59544 6520
rect 54720 6480 59544 6508
rect 54720 6468 54726 6480
rect 59538 6468 59544 6480
rect 59596 6468 59602 6520
rect 59630 6468 59636 6520
rect 59688 6508 59694 6520
rect 63770 6508 63776 6520
rect 59688 6480 63776 6508
rect 59688 6468 59694 6480
rect 63770 6468 63776 6480
rect 63828 6468 63834 6520
rect 64046 6468 64052 6520
rect 64104 6508 64110 6520
rect 64322 6508 64328 6520
rect 64104 6480 64328 6508
rect 64104 6468 64110 6480
rect 64322 6468 64328 6480
rect 64380 6468 64386 6520
rect 65320 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74980 6554
rect 65320 6480 74980 6502
rect 29546 6400 29552 6452
rect 29604 6440 29610 6452
rect 47486 6440 47492 6452
rect 29604 6412 47492 6440
rect 29604 6400 29610 6412
rect 47486 6400 47492 6412
rect 47544 6400 47550 6452
rect 49602 6400 49608 6452
rect 49660 6440 49666 6452
rect 63862 6440 63868 6452
rect 49660 6412 63868 6440
rect 49660 6400 49666 6412
rect 63862 6400 63868 6412
rect 63920 6400 63926 6452
rect 64230 6400 64236 6452
rect 64288 6440 64294 6452
rect 66438 6440 66444 6452
rect 64288 6412 66444 6440
rect 64288 6400 64294 6412
rect 66438 6400 66444 6412
rect 66496 6400 66502 6452
rect 23658 6332 23664 6384
rect 23716 6372 23722 6384
rect 32306 6372 32312 6384
rect 23716 6344 32312 6372
rect 23716 6332 23722 6344
rect 32306 6332 32312 6344
rect 32364 6332 32370 6384
rect 48130 6332 48136 6384
rect 48188 6372 48194 6384
rect 64414 6372 64420 6384
rect 48188 6344 64420 6372
rect 48188 6332 48194 6344
rect 64414 6332 64420 6344
rect 64472 6332 64478 6384
rect 65518 6332 65524 6384
rect 65576 6372 65582 6384
rect 66714 6372 66720 6384
rect 65576 6344 66720 6372
rect 65576 6332 65582 6344
rect 66714 6332 66720 6344
rect 66772 6332 66778 6384
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 34882 6304 34888 6316
rect 26200 6276 34888 6304
rect 26200 6264 26206 6276
rect 34882 6264 34888 6276
rect 34940 6264 34946 6316
rect 53926 6264 53932 6316
rect 53984 6304 53990 6316
rect 59906 6304 59912 6316
rect 53984 6276 59912 6304
rect 53984 6264 53990 6276
rect 59906 6264 59912 6276
rect 59964 6264 59970 6316
rect 59998 6264 60004 6316
rect 60056 6304 60062 6316
rect 67818 6304 67824 6316
rect 60056 6276 67824 6304
rect 60056 6264 60062 6276
rect 67818 6264 67824 6276
rect 67876 6264 67882 6316
rect 27062 6196 27068 6248
rect 27120 6236 27126 6248
rect 45646 6236 45652 6248
rect 27120 6208 45652 6236
rect 27120 6196 27126 6208
rect 45646 6196 45652 6208
rect 45704 6196 45710 6248
rect 51074 6196 51080 6248
rect 51132 6236 51138 6248
rect 55582 6236 55588 6248
rect 51132 6208 55588 6236
rect 51132 6196 51138 6208
rect 55582 6196 55588 6208
rect 55640 6196 55646 6248
rect 64322 6236 64328 6248
rect 55876 6208 64328 6236
rect 24946 6128 24952 6180
rect 25004 6168 25010 6180
rect 44910 6168 44916 6180
rect 25004 6140 44916 6168
rect 25004 6128 25010 6140
rect 44910 6128 44916 6140
rect 44968 6128 44974 6180
rect 47026 6128 47032 6180
rect 47084 6168 47090 6180
rect 55766 6168 55772 6180
rect 47084 6140 55772 6168
rect 47084 6128 47090 6140
rect 55766 6128 55772 6140
rect 55824 6128 55830 6180
rect 46290 6060 46296 6112
rect 46348 6100 46354 6112
rect 55876 6100 55904 6208
rect 64322 6196 64328 6208
rect 64380 6196 64386 6248
rect 64966 6196 64972 6248
rect 65024 6236 65030 6248
rect 66530 6236 66536 6248
rect 65024 6208 66536 6236
rect 65024 6196 65030 6208
rect 66530 6196 66536 6208
rect 66588 6196 66594 6248
rect 56042 6128 56048 6180
rect 56100 6168 56106 6180
rect 64506 6168 64512 6180
rect 56100 6140 64512 6168
rect 56100 6128 56106 6140
rect 64506 6128 64512 6140
rect 64564 6128 64570 6180
rect 46348 6072 55904 6100
rect 46348 6060 46354 6072
rect 55950 6060 55956 6112
rect 56008 6100 56014 6112
rect 63034 6100 63040 6112
rect 56008 6072 63040 6100
rect 56008 6060 56014 6072
rect 63034 6060 63040 6072
rect 63092 6060 63098 6112
rect 63126 6060 63132 6112
rect 63184 6100 63190 6112
rect 67726 6100 67732 6112
rect 63184 6072 67732 6100
rect 63184 6060 63190 6072
rect 67726 6060 67732 6072
rect 67784 6060 67790 6112
rect 1012 6010 74980 6032
rect 1012 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 74980 6010
rect 1012 5936 74980 5958
rect 23658 5856 23664 5908
rect 23716 5856 23722 5908
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 33318 5896 33324 5908
rect 24167 5868 33324 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 33318 5856 33324 5868
rect 33376 5856 33382 5908
rect 33870 5856 33876 5908
rect 33928 5896 33934 5908
rect 48958 5896 48964 5908
rect 33928 5868 48964 5896
rect 33928 5856 33934 5868
rect 48958 5856 48964 5868
rect 49016 5856 49022 5908
rect 49602 5856 49608 5908
rect 49660 5856 49666 5908
rect 51077 5899 51135 5905
rect 51077 5865 51089 5899
rect 51123 5896 51135 5899
rect 55674 5896 55680 5908
rect 51123 5868 55680 5896
rect 51123 5865 51135 5868
rect 51077 5859 51135 5865
rect 55674 5856 55680 5868
rect 55732 5856 55738 5908
rect 55766 5856 55772 5908
rect 55824 5896 55830 5908
rect 59814 5896 59820 5908
rect 55824 5868 59820 5896
rect 55824 5856 55830 5868
rect 59814 5856 59820 5868
rect 59872 5856 59878 5908
rect 59906 5856 59912 5908
rect 59964 5896 59970 5908
rect 63034 5896 63040 5908
rect 59964 5868 63040 5896
rect 59964 5856 59970 5868
rect 63034 5856 63040 5868
rect 63092 5856 63098 5908
rect 63310 5856 63316 5908
rect 63368 5896 63374 5908
rect 65426 5896 65432 5908
rect 63368 5868 65432 5896
rect 63368 5856 63374 5868
rect 65426 5856 65432 5868
rect 65484 5856 65490 5908
rect 55950 5828 55956 5840
rect 23768 5800 55956 5828
rect 23290 5720 23296 5772
rect 23348 5720 23354 5772
rect 23768 5769 23796 5800
rect 55950 5788 55956 5800
rect 56008 5788 56014 5840
rect 56137 5831 56195 5837
rect 56137 5797 56149 5831
rect 56183 5828 56195 5831
rect 56226 5828 56232 5840
rect 56183 5800 56232 5828
rect 56183 5797 56195 5800
rect 56137 5791 56195 5797
rect 56226 5788 56232 5800
rect 56284 5788 56290 5840
rect 61470 5828 61476 5840
rect 56336 5800 61476 5828
rect 23753 5763 23811 5769
rect 23753 5729 23765 5763
rect 23799 5729 23811 5763
rect 23753 5723 23811 5729
rect 24305 5763 24363 5769
rect 24305 5729 24317 5763
rect 24351 5760 24363 5763
rect 24578 5760 24584 5772
rect 24351 5732 24584 5760
rect 24351 5729 24363 5732
rect 24305 5723 24363 5729
rect 24578 5720 24584 5732
rect 24636 5720 24642 5772
rect 24673 5763 24731 5769
rect 24673 5729 24685 5763
rect 24719 5760 24731 5763
rect 32214 5760 32220 5772
rect 24719 5732 32220 5760
rect 24719 5729 24731 5732
rect 24673 5723 24731 5729
rect 32214 5720 32220 5732
rect 32272 5720 32278 5772
rect 32582 5720 32588 5772
rect 32640 5760 32646 5772
rect 48225 5763 48283 5769
rect 48225 5760 48237 5763
rect 32640 5732 48237 5760
rect 32640 5720 32646 5732
rect 48225 5729 48237 5732
rect 48271 5729 48283 5763
rect 48225 5723 48283 5729
rect 48866 5720 48872 5772
rect 48924 5720 48930 5772
rect 48958 5720 48964 5772
rect 49016 5720 49022 5772
rect 54662 5760 54668 5772
rect 49068 5732 54668 5760
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 23937 5695 23995 5701
rect 23937 5692 23949 5695
rect 23523 5664 23949 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 23937 5661 23949 5664
rect 23983 5692 23995 5695
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 23983 5664 24501 5692
rect 23983 5661 23995 5664
rect 23937 5655 23995 5661
rect 24489 5661 24501 5664
rect 24535 5661 24547 5695
rect 24489 5655 24547 5661
rect 24504 5624 24532 5655
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 24964 5624 24992 5655
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 25958 5652 25964 5704
rect 26016 5652 26022 5704
rect 26142 5652 26148 5704
rect 26200 5652 26206 5704
rect 40402 5652 40408 5704
rect 40460 5652 40466 5704
rect 41506 5652 41512 5704
rect 41564 5692 41570 5704
rect 42337 5695 42395 5701
rect 42337 5692 42349 5695
rect 41564 5664 42349 5692
rect 41564 5652 41570 5664
rect 42337 5661 42349 5664
rect 42383 5661 42395 5695
rect 42337 5655 42395 5661
rect 43806 5652 43812 5704
rect 43864 5652 43870 5704
rect 44453 5695 44511 5701
rect 44453 5661 44465 5695
rect 44499 5692 44511 5695
rect 44634 5692 44640 5704
rect 44499 5664 44640 5692
rect 44499 5661 44511 5664
rect 44453 5655 44511 5661
rect 44634 5652 44640 5664
rect 44692 5652 44698 5704
rect 44910 5652 44916 5704
rect 44968 5652 44974 5704
rect 45646 5652 45652 5704
rect 45704 5652 45710 5704
rect 46290 5652 46296 5704
rect 46348 5652 46354 5704
rect 46382 5652 46388 5704
rect 46440 5652 46446 5704
rect 47026 5652 47032 5704
rect 47084 5652 47090 5704
rect 47486 5652 47492 5704
rect 47544 5652 47550 5704
rect 49068 5692 49096 5732
rect 54662 5720 54668 5732
rect 54720 5720 54726 5772
rect 54757 5763 54815 5769
rect 54757 5729 54769 5763
rect 54803 5760 54815 5763
rect 56336 5760 56364 5800
rect 61470 5788 61476 5800
rect 61528 5788 61534 5840
rect 63862 5828 63868 5840
rect 61580 5800 63868 5828
rect 54803 5732 56364 5760
rect 54803 5729 54815 5732
rect 54757 5723 54815 5729
rect 56502 5720 56508 5772
rect 56560 5720 56566 5772
rect 57790 5720 57796 5772
rect 57848 5720 57854 5772
rect 58158 5720 58164 5772
rect 58216 5720 58222 5772
rect 58250 5720 58256 5772
rect 58308 5760 58314 5772
rect 59630 5760 59636 5772
rect 58308 5732 59636 5760
rect 58308 5720 58314 5732
rect 59630 5720 59636 5732
rect 59688 5720 59694 5772
rect 59722 5720 59728 5772
rect 59780 5720 59786 5772
rect 59814 5720 59820 5772
rect 59872 5760 59878 5772
rect 61580 5760 61608 5800
rect 63862 5788 63868 5800
rect 63920 5788 63926 5840
rect 67634 5828 67640 5840
rect 63972 5800 67640 5828
rect 59872 5732 61608 5760
rect 59872 5720 59878 5732
rect 61654 5720 61660 5772
rect 61712 5720 61718 5772
rect 62942 5720 62948 5772
rect 63000 5720 63006 5772
rect 63034 5720 63040 5772
rect 63092 5760 63098 5772
rect 63972 5760 64000 5800
rect 67634 5788 67640 5800
rect 67692 5788 67698 5840
rect 63092 5732 64000 5760
rect 63092 5720 63098 5732
rect 64046 5720 64052 5772
rect 64104 5760 64110 5772
rect 64598 5760 64604 5772
rect 64104 5732 64604 5760
rect 64104 5720 64110 5732
rect 64598 5720 64604 5732
rect 64656 5720 64662 5772
rect 65058 5720 65064 5772
rect 65116 5720 65122 5772
rect 66162 5720 66168 5772
rect 66220 5720 66226 5772
rect 68462 5720 68468 5772
rect 68520 5720 68526 5772
rect 47964 5664 49096 5692
rect 25976 5624 26004 5652
rect 24504 5596 26004 5624
rect 36998 5584 37004 5636
rect 37056 5584 37062 5636
rect 43533 5627 43591 5633
rect 43533 5593 43545 5627
rect 43579 5624 43591 5627
rect 47854 5624 47860 5636
rect 43579 5596 47860 5624
rect 43579 5593 43591 5596
rect 43533 5587 43591 5593
rect 47854 5584 47860 5596
rect 47912 5584 47918 5636
rect 25133 5559 25191 5565
rect 25133 5525 25145 5559
rect 25179 5556 25191 5559
rect 31662 5556 31668 5568
rect 25179 5528 31668 5556
rect 25179 5525 25191 5528
rect 25133 5519 25191 5525
rect 31662 5516 31668 5528
rect 31720 5516 31726 5568
rect 35713 5559 35771 5565
rect 35713 5525 35725 5559
rect 35759 5556 35771 5559
rect 35894 5556 35900 5568
rect 35759 5528 35900 5556
rect 35759 5525 35771 5528
rect 35713 5519 35771 5525
rect 35894 5516 35900 5528
rect 35952 5516 35958 5568
rect 41690 5516 41696 5568
rect 41748 5516 41754 5568
rect 45557 5559 45615 5565
rect 45557 5525 45569 5559
rect 45603 5556 45615 5559
rect 47964 5556 47992 5664
rect 50430 5652 50436 5704
rect 50488 5652 50494 5704
rect 51258 5652 51264 5704
rect 51316 5652 51322 5704
rect 51905 5695 51963 5701
rect 51905 5661 51917 5695
rect 51951 5692 51963 5695
rect 52270 5692 52276 5704
rect 51951 5664 52276 5692
rect 51951 5661 51963 5664
rect 51905 5655 51963 5661
rect 52270 5652 52276 5664
rect 52328 5652 52334 5704
rect 52638 5652 52644 5704
rect 52696 5652 52702 5704
rect 53374 5652 53380 5704
rect 53432 5652 53438 5704
rect 53926 5652 53932 5704
rect 53984 5692 53990 5704
rect 54021 5695 54079 5701
rect 54021 5692 54033 5695
rect 53984 5664 54033 5692
rect 53984 5652 53990 5664
rect 54021 5661 54033 5664
rect 54067 5661 54079 5695
rect 54021 5655 54079 5661
rect 54205 5695 54263 5701
rect 54205 5661 54217 5695
rect 54251 5692 54263 5695
rect 54570 5692 54576 5704
rect 54251 5664 54576 5692
rect 54251 5661 54263 5664
rect 54205 5655 54263 5661
rect 54570 5652 54576 5664
rect 54628 5652 54634 5704
rect 55306 5652 55312 5704
rect 55364 5652 55370 5704
rect 55861 5695 55919 5701
rect 55861 5661 55873 5695
rect 55907 5692 55919 5695
rect 56134 5692 56140 5704
rect 55907 5664 56140 5692
rect 55907 5661 55919 5664
rect 55861 5655 55919 5661
rect 56134 5652 56140 5664
rect 56192 5652 56198 5704
rect 56318 5652 56324 5704
rect 56376 5692 56382 5704
rect 57977 5695 58035 5701
rect 57977 5692 57989 5695
rect 56376 5664 57989 5692
rect 56376 5652 56382 5664
rect 57977 5661 57989 5664
rect 58023 5692 58035 5695
rect 59541 5695 59599 5701
rect 59541 5692 59553 5695
rect 58023 5664 59553 5692
rect 58023 5661 58035 5664
rect 57977 5655 58035 5661
rect 59541 5661 59553 5664
rect 59587 5692 59599 5695
rect 61102 5692 61108 5704
rect 59587 5664 61108 5692
rect 59587 5661 59599 5664
rect 59541 5655 59599 5661
rect 61102 5652 61108 5664
rect 61160 5692 61166 5704
rect 61473 5695 61531 5701
rect 61473 5692 61485 5695
rect 61160 5664 61485 5692
rect 61160 5652 61166 5664
rect 61473 5661 61485 5664
rect 61519 5692 61531 5695
rect 63129 5695 63187 5701
rect 63129 5692 63141 5695
rect 61519 5664 63141 5692
rect 61519 5661 61531 5664
rect 61473 5655 61531 5661
rect 63129 5661 63141 5664
rect 63175 5692 63187 5695
rect 64877 5695 64935 5701
rect 64877 5692 64889 5695
rect 63175 5664 64889 5692
rect 63175 5661 63187 5664
rect 63129 5655 63187 5661
rect 64877 5661 64889 5664
rect 64923 5692 64935 5695
rect 66349 5695 66407 5701
rect 66349 5692 66361 5695
rect 64923 5664 66361 5692
rect 64923 5661 64935 5664
rect 64877 5655 64935 5661
rect 66349 5661 66361 5664
rect 66395 5692 66407 5695
rect 68281 5695 68339 5701
rect 68281 5692 68293 5695
rect 66395 5664 68293 5692
rect 66395 5661 66407 5664
rect 66349 5655 66407 5661
rect 68281 5661 68293 5664
rect 68327 5661 68339 5695
rect 68281 5655 68339 5661
rect 48038 5584 48044 5636
rect 48096 5624 48102 5636
rect 61010 5624 61016 5636
rect 48096 5596 61016 5624
rect 48096 5584 48102 5596
rect 61010 5584 61016 5596
rect 61068 5584 61074 5636
rect 64046 5624 64052 5636
rect 61120 5596 64052 5624
rect 45603 5528 47992 5556
rect 45603 5525 45615 5528
rect 45557 5519 45615 5525
rect 48130 5516 48136 5568
rect 48188 5516 48194 5568
rect 53285 5559 53343 5565
rect 53285 5525 53297 5559
rect 53331 5556 53343 5559
rect 58250 5556 58256 5568
rect 53331 5528 58256 5556
rect 53331 5525 53343 5528
rect 53285 5519 53343 5525
rect 58250 5516 58256 5528
rect 58308 5516 58314 5568
rect 59357 5559 59415 5565
rect 59357 5525 59369 5559
rect 59403 5556 59415 5559
rect 59446 5556 59452 5568
rect 59403 5528 59452 5556
rect 59403 5525 59415 5528
rect 59357 5519 59415 5525
rect 59446 5516 59452 5528
rect 59504 5516 59510 5568
rect 59538 5516 59544 5568
rect 59596 5556 59602 5568
rect 61120 5556 61148 5596
rect 64046 5584 64052 5596
rect 64104 5584 64110 5636
rect 68830 5624 68836 5636
rect 64616 5596 68836 5624
rect 59596 5528 61148 5556
rect 59596 5516 59602 5528
rect 61194 5516 61200 5568
rect 61252 5556 61258 5568
rect 61289 5559 61347 5565
rect 61289 5556 61301 5559
rect 61252 5528 61301 5556
rect 61252 5516 61258 5528
rect 61289 5525 61301 5528
rect 61335 5525 61347 5559
rect 61289 5519 61347 5525
rect 61470 5516 61476 5568
rect 61528 5556 61534 5568
rect 63126 5556 63132 5568
rect 61528 5528 63132 5556
rect 61528 5516 61534 5528
rect 63126 5516 63132 5528
rect 63184 5516 63190 5568
rect 63218 5516 63224 5568
rect 63276 5556 63282 5568
rect 63313 5559 63371 5565
rect 63313 5556 63325 5559
rect 63276 5528 63325 5556
rect 63276 5516 63282 5528
rect 63313 5525 63325 5528
rect 63359 5525 63371 5559
rect 63313 5519 63371 5525
rect 63402 5516 63408 5568
rect 63460 5556 63466 5568
rect 64616 5556 64644 5596
rect 68830 5584 68836 5596
rect 68888 5584 68894 5636
rect 63460 5528 64644 5556
rect 64693 5559 64751 5565
rect 63460 5516 63466 5528
rect 64693 5525 64705 5559
rect 64739 5556 64751 5559
rect 64782 5556 64788 5568
rect 64739 5528 64788 5556
rect 64739 5525 64751 5528
rect 64693 5519 64751 5525
rect 64782 5516 64788 5528
rect 64840 5516 64846 5568
rect 66438 5516 66444 5568
rect 66496 5556 66502 5568
rect 66533 5559 66591 5565
rect 66533 5556 66545 5559
rect 66496 5528 66545 5556
rect 66496 5516 66502 5528
rect 66533 5525 66545 5528
rect 66579 5525 66591 5559
rect 66533 5519 66591 5525
rect 68094 5516 68100 5568
rect 68152 5516 68158 5568
rect 1012 5466 74980 5488
rect 1012 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74980 5466
rect 1012 5392 74980 5414
rect 25958 5352 25964 5364
rect 25700 5324 25964 5352
rect 24412 5256 25544 5284
rect 23934 5176 23940 5228
rect 23992 5216 23998 5228
rect 24412 5225 24440 5256
rect 24397 5219 24455 5225
rect 24397 5216 24409 5219
rect 23992 5188 24409 5216
rect 23992 5176 23998 5188
rect 24397 5185 24409 5188
rect 24443 5185 24455 5219
rect 24397 5179 24455 5185
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5148 24271 5151
rect 24578 5148 24584 5160
rect 24259 5120 24584 5148
rect 24259 5117 24271 5120
rect 24213 5111 24271 5117
rect 24578 5108 24584 5120
rect 24636 5108 24642 5160
rect 25406 5108 25412 5160
rect 25464 5108 25470 5160
rect 25516 5148 25544 5256
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5216 25651 5219
rect 25700 5216 25728 5324
rect 25958 5312 25964 5324
rect 26016 5352 26022 5364
rect 27798 5352 27804 5364
rect 26016 5324 27804 5352
rect 26016 5312 26022 5324
rect 27798 5312 27804 5324
rect 27856 5312 27862 5364
rect 27893 5355 27951 5361
rect 27893 5321 27905 5355
rect 27939 5352 27951 5355
rect 36814 5352 36820 5364
rect 27939 5324 36820 5352
rect 27939 5321 27951 5324
rect 27893 5315 27951 5321
rect 36814 5312 36820 5324
rect 36872 5312 36878 5364
rect 41046 5312 41052 5364
rect 41104 5312 41110 5364
rect 41138 5312 41144 5364
rect 41196 5352 41202 5364
rect 54754 5352 54760 5364
rect 41196 5324 54760 5352
rect 41196 5312 41202 5324
rect 54754 5312 54760 5324
rect 54812 5312 54818 5364
rect 60642 5352 60648 5364
rect 54864 5324 60648 5352
rect 27614 5284 27620 5296
rect 27264 5256 27620 5284
rect 27264 5225 27292 5256
rect 27614 5244 27620 5256
rect 27672 5284 27678 5296
rect 27672 5256 27936 5284
rect 27672 5244 27678 5256
rect 26053 5219 26111 5225
rect 26053 5216 26065 5219
rect 25639 5188 25728 5216
rect 25792 5188 26065 5216
rect 25639 5185 25651 5188
rect 25593 5179 25651 5185
rect 25792 5148 25820 5188
rect 26053 5185 26065 5188
rect 26099 5216 26111 5219
rect 26513 5219 26571 5225
rect 27249 5222 27307 5225
rect 26513 5216 26525 5219
rect 26099 5188 26525 5216
rect 26099 5185 26111 5188
rect 26053 5179 26111 5185
rect 26513 5185 26525 5188
rect 26559 5216 26571 5219
rect 27080 5219 27307 5222
rect 26559 5214 27016 5216
rect 27080 5214 27261 5219
rect 26559 5194 27261 5214
rect 26559 5188 27108 5194
rect 26559 5185 26571 5188
rect 26988 5186 27108 5188
rect 26513 5179 26571 5185
rect 27249 5185 27261 5194
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27430 5176 27436 5228
rect 27488 5216 27494 5228
rect 27709 5219 27767 5225
rect 27488 5188 27660 5216
rect 27488 5176 27494 5188
rect 25516 5120 25820 5148
rect 25869 5151 25927 5157
rect 25869 5117 25881 5151
rect 25915 5117 25927 5151
rect 25869 5111 25927 5117
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 24673 5083 24731 5089
rect 24673 5080 24685 5083
rect 23532 5052 24685 5080
rect 23532 5040 23538 5052
rect 24673 5049 24685 5052
rect 24719 5049 24731 5083
rect 24673 5043 24731 5049
rect 25774 5040 25780 5092
rect 25832 5040 25838 5092
rect 25884 5080 25912 5111
rect 26326 5108 26332 5160
rect 26384 5108 26390 5160
rect 27065 5151 27123 5157
rect 27065 5117 27077 5151
rect 27111 5148 27123 5151
rect 27154 5148 27160 5160
rect 27111 5120 27160 5148
rect 27111 5117 27123 5120
rect 27065 5111 27123 5117
rect 27154 5108 27160 5120
rect 27212 5108 27218 5160
rect 27522 5108 27528 5160
rect 27580 5108 27586 5160
rect 27632 5148 27660 5188
rect 27709 5185 27721 5219
rect 27755 5216 27767 5219
rect 27798 5216 27804 5228
rect 27755 5188 27804 5216
rect 27755 5185 27767 5188
rect 27709 5179 27767 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 27908 5216 27936 5256
rect 28074 5244 28080 5296
rect 28132 5284 28138 5296
rect 31202 5284 31208 5296
rect 28132 5256 31208 5284
rect 28132 5244 28138 5256
rect 31202 5244 31208 5256
rect 31260 5244 31266 5296
rect 54662 5284 54668 5296
rect 31312 5256 41092 5284
rect 28261 5219 28319 5225
rect 28261 5216 28273 5219
rect 27908 5188 28273 5216
rect 28261 5185 28273 5188
rect 28307 5216 28319 5219
rect 28905 5219 28963 5225
rect 28905 5216 28917 5219
rect 28307 5188 28917 5216
rect 28307 5185 28319 5188
rect 28261 5179 28319 5185
rect 28905 5185 28917 5188
rect 28951 5216 28963 5219
rect 29549 5219 29607 5225
rect 29549 5216 29561 5219
rect 28951 5188 29561 5216
rect 28951 5185 28963 5188
rect 28905 5179 28963 5185
rect 29549 5185 29561 5188
rect 29595 5216 29607 5219
rect 30101 5219 30159 5225
rect 30101 5216 30113 5219
rect 29595 5188 30113 5216
rect 29595 5185 29607 5188
rect 29549 5179 29607 5185
rect 30101 5185 30113 5188
rect 30147 5185 30159 5219
rect 30101 5179 30159 5185
rect 27632 5120 28396 5148
rect 27246 5080 27252 5092
rect 25884 5052 27252 5080
rect 27246 5040 27252 5052
rect 27304 5040 27310 5092
rect 27433 5083 27491 5089
rect 27433 5049 27445 5083
rect 27479 5080 27491 5083
rect 28258 5080 28264 5092
rect 27479 5052 28264 5080
rect 27479 5049 27491 5052
rect 27433 5043 27491 5049
rect 28258 5040 28264 5052
rect 28316 5040 28322 5092
rect 28368 5080 28396 5120
rect 28442 5108 28448 5160
rect 28500 5108 28506 5160
rect 29086 5108 29092 5160
rect 29144 5108 29150 5160
rect 29730 5108 29736 5160
rect 29788 5108 29794 5160
rect 30116 5148 30144 5179
rect 30282 5176 30288 5228
rect 30340 5176 30346 5228
rect 30653 5219 30711 5225
rect 30653 5185 30665 5219
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 30668 5148 30696 5179
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 30116 5120 30696 5148
rect 31312 5080 31340 5256
rect 31386 5176 31392 5228
rect 31444 5216 31450 5228
rect 40954 5216 40960 5228
rect 31444 5188 40960 5216
rect 31444 5176 31450 5188
rect 40954 5176 40960 5188
rect 41012 5176 41018 5228
rect 41064 5216 41092 5256
rect 41386 5256 54668 5284
rect 41386 5216 41414 5256
rect 54662 5244 54668 5256
rect 54720 5244 54726 5296
rect 41064 5188 41414 5216
rect 41690 5176 41696 5228
rect 41748 5216 41754 5228
rect 42981 5219 43039 5225
rect 42981 5216 42993 5219
rect 41748 5188 42993 5216
rect 41748 5176 41754 5188
rect 42981 5185 42993 5188
rect 43027 5185 43039 5219
rect 42981 5179 43039 5185
rect 44177 5219 44235 5225
rect 44177 5185 44189 5219
rect 44223 5216 44235 5219
rect 44223 5188 46152 5216
rect 44223 5185 44235 5188
rect 44177 5179 44235 5185
rect 40402 5108 40408 5160
rect 40460 5108 40466 5160
rect 41509 5151 41567 5157
rect 41509 5148 41521 5151
rect 41386 5120 41521 5148
rect 28368 5052 31340 5080
rect 40586 5040 40592 5092
rect 40644 5080 40650 5092
rect 41386 5080 41414 5120
rect 41509 5117 41521 5120
rect 41555 5117 41567 5151
rect 41509 5111 41567 5117
rect 42153 5151 42211 5157
rect 42153 5117 42165 5151
rect 42199 5148 42211 5151
rect 42702 5148 42708 5160
rect 42199 5120 42708 5148
rect 42199 5117 42211 5120
rect 42153 5111 42211 5117
rect 42702 5108 42708 5120
rect 42760 5108 42766 5160
rect 44545 5151 44603 5157
rect 44545 5117 44557 5151
rect 44591 5117 44603 5151
rect 45373 5151 45431 5157
rect 45373 5148 45385 5151
rect 44545 5111 44603 5117
rect 44744 5120 45385 5148
rect 40644 5052 41414 5080
rect 44560 5080 44588 5111
rect 44634 5080 44640 5092
rect 44560 5052 44640 5080
rect 40644 5040 40650 5052
rect 44634 5040 44640 5052
rect 44692 5040 44698 5092
rect 24581 5015 24639 5021
rect 24581 4981 24593 5015
rect 24627 5012 24639 5015
rect 26142 5012 26148 5024
rect 24627 4984 26148 5012
rect 24627 4981 24639 4984
rect 24581 4975 24639 4981
rect 26142 4972 26148 4984
rect 26200 4972 26206 5024
rect 26234 4972 26240 5024
rect 26292 4972 26298 5024
rect 26694 4972 26700 5024
rect 26752 4972 26758 5024
rect 28077 5015 28135 5021
rect 28077 4981 28089 5015
rect 28123 5012 28135 5015
rect 28534 5012 28540 5024
rect 28123 4984 28540 5012
rect 28123 4981 28135 4984
rect 28077 4975 28135 4981
rect 28534 4972 28540 4984
rect 28592 4972 28598 5024
rect 28718 4972 28724 5024
rect 28776 4972 28782 5024
rect 29362 4972 29368 5024
rect 29420 4972 29426 5024
rect 29454 4972 29460 5024
rect 29512 5012 29518 5024
rect 29917 5015 29975 5021
rect 29917 5012 29929 5015
rect 29512 4984 29929 5012
rect 29512 4972 29518 4984
rect 29917 4981 29929 4984
rect 29963 4981 29975 5015
rect 29917 4975 29975 4981
rect 30466 4972 30472 5024
rect 30524 4972 30530 5024
rect 33042 4972 33048 5024
rect 33100 5012 33106 5024
rect 44744 5012 44772 5120
rect 45373 5117 45385 5120
rect 45419 5117 45431 5151
rect 46124 5148 46152 5188
rect 46198 5176 46204 5228
rect 46256 5176 46262 5228
rect 46290 5176 46296 5228
rect 46348 5176 46354 5228
rect 47213 5219 47271 5225
rect 46492 5188 47164 5216
rect 46492 5148 46520 5188
rect 46124 5120 46520 5148
rect 45373 5111 45431 5117
rect 46566 5108 46572 5160
rect 46624 5108 46630 5160
rect 47136 5148 47164 5188
rect 47213 5185 47225 5219
rect 47259 5216 47271 5219
rect 53006 5216 53012 5228
rect 47259 5188 53012 5216
rect 47259 5185 47271 5188
rect 47213 5179 47271 5185
rect 53006 5176 53012 5188
rect 53064 5176 53070 5228
rect 54864 5225 54892 5324
rect 60642 5312 60648 5324
rect 60700 5312 60706 5364
rect 65886 5352 65892 5364
rect 60844 5324 65892 5352
rect 55030 5244 55036 5296
rect 55088 5284 55094 5296
rect 60844 5284 60872 5324
rect 65886 5312 65892 5324
rect 65944 5312 65950 5364
rect 65334 5284 65340 5296
rect 55088 5256 60872 5284
rect 60936 5256 65340 5284
rect 55088 5244 55094 5256
rect 53101 5219 53159 5225
rect 53101 5185 53113 5219
rect 53147 5216 53159 5219
rect 54757 5219 54815 5225
rect 54757 5216 54769 5219
rect 53147 5188 54769 5216
rect 53147 5185 53159 5188
rect 53101 5179 53159 5185
rect 54757 5185 54769 5188
rect 54803 5185 54815 5219
rect 54757 5179 54815 5185
rect 54849 5219 54907 5225
rect 54849 5185 54861 5219
rect 54895 5185 54907 5219
rect 56318 5216 56324 5228
rect 54849 5179 54907 5185
rect 55048 5188 56324 5216
rect 47136 5120 47348 5148
rect 45097 5083 45155 5089
rect 45097 5049 45109 5083
rect 45143 5080 45155 5083
rect 47210 5080 47216 5092
rect 45143 5052 47216 5080
rect 45143 5049 45155 5052
rect 45097 5043 45155 5049
rect 47210 5040 47216 5052
rect 47268 5040 47274 5092
rect 33100 4984 44772 5012
rect 33100 4972 33106 4984
rect 46014 4972 46020 5024
rect 46072 4972 46078 5024
rect 46477 5015 46535 5021
rect 46477 4981 46489 5015
rect 46523 5012 46535 5015
rect 47118 5012 47124 5024
rect 46523 4984 47124 5012
rect 46523 4981 46535 4984
rect 46477 4975 46535 4981
rect 47118 4972 47124 4984
rect 47176 4972 47182 5024
rect 47320 5012 47348 5120
rect 47486 5108 47492 5160
rect 47544 5108 47550 5160
rect 48133 5151 48191 5157
rect 48133 5117 48145 5151
rect 48179 5148 48191 5151
rect 48222 5148 48228 5160
rect 48179 5120 48228 5148
rect 48179 5117 48191 5120
rect 48133 5111 48191 5117
rect 48222 5108 48228 5120
rect 48280 5108 48286 5160
rect 49142 5108 49148 5160
rect 49200 5108 49206 5160
rect 49789 5151 49847 5157
rect 49789 5117 49801 5151
rect 49835 5148 49847 5151
rect 50982 5148 50988 5160
rect 49835 5120 50988 5148
rect 49835 5117 49847 5120
rect 49789 5111 49847 5117
rect 50982 5108 50988 5120
rect 51040 5108 51046 5160
rect 53282 5108 53288 5160
rect 53340 5108 53346 5160
rect 54772 5148 54800 5179
rect 55048 5148 55076 5188
rect 56318 5176 56324 5188
rect 56376 5176 56382 5228
rect 56410 5176 56416 5228
rect 56468 5216 56474 5228
rect 56468 5214 60780 5216
rect 60936 5214 60964 5256
rect 65334 5244 65340 5256
rect 65392 5244 65398 5296
rect 69658 5244 69664 5296
rect 69716 5284 69722 5296
rect 69716 5256 73568 5284
rect 69716 5244 69722 5256
rect 56468 5188 60964 5214
rect 56468 5176 56474 5188
rect 60752 5186 60964 5188
rect 61286 5176 61292 5228
rect 61344 5216 61350 5228
rect 73540 5225 73568 5256
rect 70213 5219 70271 5225
rect 70213 5216 70225 5219
rect 61344 5188 70225 5216
rect 61344 5176 61350 5188
rect 70213 5185 70225 5188
rect 70259 5216 70271 5219
rect 71685 5219 71743 5225
rect 71685 5216 71697 5219
rect 70259 5188 71697 5216
rect 70259 5185 70271 5188
rect 70213 5179 70271 5185
rect 71685 5185 71697 5188
rect 71731 5216 71743 5219
rect 73433 5219 73491 5225
rect 73433 5216 73445 5219
rect 71731 5188 73445 5216
rect 71731 5185 71743 5188
rect 71685 5179 71743 5185
rect 73433 5185 73445 5188
rect 73479 5185 73491 5219
rect 73433 5179 73491 5185
rect 73525 5219 73583 5225
rect 73525 5185 73537 5219
rect 73571 5185 73583 5219
rect 73525 5179 73583 5185
rect 54772 5120 55076 5148
rect 55122 5108 55128 5160
rect 55180 5148 55186 5160
rect 65610 5148 65616 5160
rect 55180 5120 65616 5148
rect 55180 5108 55186 5120
rect 65610 5108 65616 5120
rect 65668 5108 65674 5160
rect 69934 5108 69940 5160
rect 69992 5148 69998 5160
rect 70397 5151 70455 5157
rect 70397 5148 70409 5151
rect 69992 5120 70409 5148
rect 69992 5108 69998 5120
rect 70397 5117 70409 5120
rect 70443 5117 70455 5151
rect 70397 5111 70455 5117
rect 71869 5151 71927 5157
rect 71869 5117 71881 5151
rect 71915 5117 71927 5151
rect 71869 5111 71927 5117
rect 47394 5040 47400 5092
rect 47452 5080 47458 5092
rect 47452 5052 55904 5080
rect 47452 5040 47458 5052
rect 49510 5012 49516 5024
rect 47320 4984 49516 5012
rect 49510 4972 49516 4984
rect 49568 4972 49574 5024
rect 52914 4972 52920 5024
rect 52972 4972 52978 5024
rect 54573 5015 54631 5021
rect 54573 4981 54585 5015
rect 54619 5012 54631 5015
rect 54662 5012 54668 5024
rect 54619 4984 54668 5012
rect 54619 4981 54631 4984
rect 54573 4975 54631 4981
rect 54662 4972 54668 4984
rect 54720 4972 54726 5024
rect 55876 5012 55904 5052
rect 55950 5040 55956 5092
rect 56008 5080 56014 5092
rect 66070 5080 66076 5092
rect 56008 5052 66076 5080
rect 56008 5040 56014 5052
rect 66070 5040 66076 5052
rect 66128 5040 66134 5092
rect 69750 5040 69756 5092
rect 69808 5080 69814 5092
rect 71884 5080 71912 5111
rect 69808 5052 71912 5080
rect 69808 5040 69814 5052
rect 68186 5012 68192 5024
rect 55876 4984 68192 5012
rect 68186 4972 68192 4984
rect 68244 4972 68250 5024
rect 69842 4972 69848 5024
rect 69900 5012 69906 5024
rect 70029 5015 70087 5021
rect 70029 5012 70041 5015
rect 69900 4984 70041 5012
rect 69900 4972 69906 4984
rect 70029 4981 70041 4984
rect 70075 4981 70087 5015
rect 70029 4975 70087 4981
rect 71406 4972 71412 5024
rect 71464 5012 71470 5024
rect 71501 5015 71559 5021
rect 71501 5012 71513 5015
rect 71464 4984 71513 5012
rect 71464 4972 71470 4984
rect 71501 4981 71513 4984
rect 71547 4981 71559 5015
rect 71501 4975 71559 4981
rect 73246 4972 73252 5024
rect 73304 4972 73310 5024
rect 1012 4922 74980 4944
rect 1012 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 74980 4922
rect 1012 4848 74980 4870
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 30006 4808 30012 4820
rect 26292 4780 30012 4808
rect 26292 4768 26298 4780
rect 30006 4768 30012 4780
rect 30064 4768 30070 4820
rect 31018 4768 31024 4820
rect 31076 4808 31082 4820
rect 40586 4808 40592 4820
rect 31076 4780 40592 4808
rect 31076 4768 31082 4780
rect 40586 4768 40592 4780
rect 40644 4768 40650 4820
rect 44726 4808 44732 4820
rect 44560 4780 44732 4808
rect 25406 4700 25412 4752
rect 25464 4740 25470 4752
rect 25464 4712 34008 4740
rect 25464 4700 25470 4712
rect 24578 4632 24584 4684
rect 24636 4672 24642 4684
rect 31386 4672 31392 4684
rect 24636 4644 31392 4672
rect 24636 4632 24642 4644
rect 31386 4632 31392 4644
rect 31444 4632 31450 4684
rect 33980 4672 34008 4712
rect 35066 4700 35072 4752
rect 35124 4740 35130 4752
rect 41690 4740 41696 4752
rect 35124 4712 41696 4740
rect 35124 4700 35130 4712
rect 41690 4700 41696 4712
rect 41748 4700 41754 4752
rect 43346 4672 43352 4684
rect 33980 4644 43352 4672
rect 43346 4632 43352 4644
rect 43404 4632 43410 4684
rect 44085 4675 44143 4681
rect 44085 4641 44097 4675
rect 44131 4672 44143 4675
rect 44560 4672 44588 4780
rect 44726 4768 44732 4780
rect 44784 4768 44790 4820
rect 46014 4768 46020 4820
rect 46072 4808 46078 4820
rect 60090 4808 60096 4820
rect 46072 4780 60096 4808
rect 46072 4768 46078 4780
rect 60090 4768 60096 4780
rect 60148 4768 60154 4820
rect 61102 4768 61108 4820
rect 61160 4768 61166 4820
rect 45094 4700 45100 4752
rect 45152 4740 45158 4752
rect 45152 4712 49372 4740
rect 45152 4700 45158 4712
rect 44131 4644 44588 4672
rect 44131 4641 44143 4644
rect 44085 4635 44143 4641
rect 44726 4632 44732 4684
rect 44784 4672 44790 4684
rect 48958 4672 48964 4684
rect 44784 4644 48964 4672
rect 44784 4632 44790 4644
rect 48958 4632 48964 4644
rect 49016 4632 49022 4684
rect 27614 4564 27620 4616
rect 27672 4604 27678 4616
rect 33778 4604 33784 4616
rect 27672 4576 33784 4604
rect 27672 4564 27678 4576
rect 33778 4564 33784 4576
rect 33836 4564 33842 4616
rect 33962 4564 33968 4616
rect 34020 4564 34026 4616
rect 34054 4564 34060 4616
rect 34112 4604 34118 4616
rect 34241 4607 34299 4613
rect 34241 4604 34253 4607
rect 34112 4576 34253 4604
rect 34112 4564 34118 4576
rect 34241 4573 34253 4576
rect 34287 4573 34299 4607
rect 34241 4567 34299 4573
rect 41230 4564 41236 4616
rect 41288 4564 41294 4616
rect 41690 4564 41696 4616
rect 41748 4604 41754 4616
rect 41969 4607 42027 4613
rect 41969 4604 41981 4607
rect 41748 4576 41981 4604
rect 41748 4564 41754 4576
rect 41969 4573 41981 4576
rect 42015 4573 42027 4607
rect 41969 4567 42027 4573
rect 43441 4607 43499 4613
rect 43441 4573 43453 4607
rect 43487 4604 43499 4607
rect 43530 4604 43536 4616
rect 43487 4576 43536 4604
rect 43487 4573 43499 4576
rect 43441 4567 43499 4573
rect 43530 4564 43536 4576
rect 43588 4564 43594 4616
rect 44269 4607 44327 4613
rect 44269 4573 44281 4607
rect 44315 4604 44327 4607
rect 46290 4604 46296 4616
rect 44315 4576 46296 4604
rect 44315 4573 44327 4576
rect 44269 4567 44327 4573
rect 26694 4496 26700 4548
rect 26752 4536 26758 4548
rect 29270 4536 29276 4548
rect 26752 4508 29276 4536
rect 26752 4496 26758 4508
rect 29270 4496 29276 4508
rect 29328 4496 29334 4548
rect 29730 4496 29736 4548
rect 29788 4536 29794 4548
rect 34698 4536 34704 4548
rect 29788 4508 34704 4536
rect 29788 4496 29794 4508
rect 34698 4496 34704 4508
rect 34756 4536 34762 4548
rect 44284 4536 44312 4567
rect 46290 4564 46296 4576
rect 46348 4604 46354 4616
rect 46658 4614 46664 4616
rect 46584 4604 46664 4614
rect 46348 4586 46664 4604
rect 46348 4576 46612 4586
rect 46348 4564 46354 4576
rect 46658 4564 46664 4586
rect 46716 4564 46722 4616
rect 46750 4564 46756 4616
rect 46808 4564 46814 4616
rect 46842 4564 46848 4616
rect 46900 4564 46906 4616
rect 34756 4508 44312 4536
rect 34756 4496 34762 4508
rect 46934 4496 46940 4548
rect 46992 4536 46998 4548
rect 49344 4536 49372 4712
rect 53006 4700 53012 4752
rect 53064 4740 53070 4752
rect 60366 4740 60372 4752
rect 53064 4712 60372 4740
rect 53064 4700 53070 4712
rect 60366 4700 60372 4712
rect 60424 4700 60430 4752
rect 62666 4740 62672 4752
rect 61212 4712 62672 4740
rect 61212 4672 61240 4712
rect 62666 4700 62672 4712
rect 62724 4700 62730 4752
rect 61120 4644 61240 4672
rect 49418 4564 49424 4616
rect 49476 4604 49482 4616
rect 61120 4604 61148 4644
rect 61378 4632 61384 4684
rect 61436 4672 61442 4684
rect 69014 4672 69020 4684
rect 61436 4644 69020 4672
rect 61436 4632 61442 4644
rect 69014 4632 69020 4644
rect 69072 4632 69078 4684
rect 49476 4576 61148 4604
rect 61197 4607 61255 4613
rect 49476 4564 49482 4576
rect 61197 4573 61209 4607
rect 61243 4604 61255 4607
rect 61286 4604 61292 4616
rect 61243 4576 61292 4604
rect 61243 4573 61255 4576
rect 61197 4567 61255 4573
rect 61286 4564 61292 4576
rect 61344 4564 61350 4616
rect 62666 4564 62672 4616
rect 62724 4604 62730 4616
rect 67910 4604 67916 4616
rect 62724 4576 67916 4604
rect 62724 4564 62730 4576
rect 67910 4564 67916 4576
rect 67968 4564 67974 4616
rect 60734 4536 60740 4548
rect 46992 4508 49188 4536
rect 49344 4508 60740 4536
rect 46992 4496 46998 4508
rect 26142 4428 26148 4480
rect 26200 4468 26206 4480
rect 29638 4468 29644 4480
rect 26200 4440 29644 4468
rect 26200 4428 26206 4440
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 33778 4428 33784 4480
rect 33836 4468 33842 4480
rect 34790 4468 34796 4480
rect 33836 4440 34796 4468
rect 33836 4428 33842 4440
rect 34790 4428 34796 4440
rect 34848 4468 34854 4480
rect 35710 4468 35716 4480
rect 34848 4440 35716 4468
rect 34848 4428 34854 4440
rect 35710 4428 35716 4440
rect 35768 4428 35774 4480
rect 41877 4471 41935 4477
rect 41877 4437 41889 4471
rect 41923 4468 41935 4471
rect 42518 4468 42524 4480
rect 41923 4440 42524 4468
rect 41923 4437 41935 4440
rect 41877 4431 41935 4437
rect 42518 4428 42524 4440
rect 42576 4428 42582 4480
rect 42610 4428 42616 4480
rect 42668 4428 42674 4480
rect 43990 4428 43996 4480
rect 44048 4428 44054 4480
rect 44453 4471 44511 4477
rect 44453 4437 44465 4471
rect 44499 4468 44511 4471
rect 45922 4468 45928 4480
rect 44499 4440 45928 4468
rect 44499 4437 44511 4440
rect 44453 4431 44511 4437
rect 45922 4428 45928 4440
rect 45980 4428 45986 4480
rect 47029 4471 47087 4477
rect 47029 4437 47041 4471
rect 47075 4468 47087 4471
rect 49050 4468 49056 4480
rect 47075 4440 49056 4468
rect 47075 4437 47087 4440
rect 47029 4431 47087 4437
rect 49050 4428 49056 4440
rect 49108 4428 49114 4480
rect 49160 4468 49188 4508
rect 60734 4496 60740 4508
rect 60792 4496 60798 4548
rect 62758 4496 62764 4548
rect 62816 4536 62822 4548
rect 68646 4536 68652 4548
rect 62816 4508 68652 4536
rect 62816 4496 62822 4508
rect 68646 4496 68652 4508
rect 68704 4496 68710 4548
rect 60826 4468 60832 4480
rect 49160 4440 60832 4468
rect 60826 4428 60832 4440
rect 60884 4428 60890 4480
rect 61010 4428 61016 4480
rect 61068 4468 61074 4480
rect 68554 4468 68560 4480
rect 61068 4440 68560 4468
rect 61068 4428 61074 4440
rect 68554 4428 68560 4440
rect 68612 4428 68618 4480
rect 1012 4378 74980 4400
rect 1012 4326 4210 4378
rect 4262 4326 4274 4378
rect 4326 4326 4338 4378
rect 4390 4326 4402 4378
rect 4454 4326 4466 4378
rect 4518 4326 14210 4378
rect 14262 4326 14274 4378
rect 14326 4326 14338 4378
rect 14390 4326 14402 4378
rect 14454 4326 14466 4378
rect 14518 4326 24210 4378
rect 24262 4326 24274 4378
rect 24326 4326 24338 4378
rect 24390 4326 24402 4378
rect 24454 4326 24466 4378
rect 24518 4326 34210 4378
rect 34262 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 44210 4378
rect 44262 4326 44274 4378
rect 44326 4326 44338 4378
rect 44390 4326 44402 4378
rect 44454 4326 44466 4378
rect 44518 4326 54210 4378
rect 54262 4326 54274 4378
rect 54326 4326 54338 4378
rect 54390 4326 54402 4378
rect 54454 4326 54466 4378
rect 54518 4326 64210 4378
rect 64262 4326 64274 4378
rect 64326 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 74210 4378
rect 74262 4326 74274 4378
rect 74326 4326 74338 4378
rect 74390 4326 74402 4378
rect 74454 4326 74466 4378
rect 74518 4326 74980 4378
rect 1012 4304 74980 4326
rect 26326 4224 26332 4276
rect 26384 4264 26390 4276
rect 63494 4264 63500 4276
rect 26384 4236 63500 4264
rect 26384 4224 26390 4236
rect 63494 4224 63500 4236
rect 63552 4224 63558 4276
rect 33042 4196 33048 4208
rect 19628 4168 20392 4196
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 19628 4128 19656 4168
rect 19116 4100 19656 4128
rect 19705 4131 19763 4137
rect 19116 4088 19122 4100
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 20254 4128 20260 4140
rect 19751 4100 20260 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20364 4128 20392 4168
rect 27540 4168 29960 4196
rect 27540 4128 27568 4168
rect 20364 4100 27568 4128
rect 27614 4088 27620 4140
rect 27672 4088 27678 4140
rect 29932 4128 29960 4168
rect 31726 4168 33048 4196
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 27724 4100 29868 4128
rect 29932 4100 30849 4128
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 27724 4060 27752 4100
rect 19567 4032 27752 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 29730 4020 29736 4072
rect 29788 4020 29794 4072
rect 29840 4060 29868 4100
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 31386 4088 31392 4140
rect 31444 4128 31450 4140
rect 31726 4128 31754 4168
rect 33042 4156 33048 4168
rect 33100 4156 33106 4208
rect 34624 4168 35020 4196
rect 31444 4100 31754 4128
rect 31444 4088 31450 4100
rect 33778 4088 33784 4140
rect 33836 4128 33842 4140
rect 34624 4128 34652 4168
rect 33836 4100 34652 4128
rect 33836 4088 33842 4100
rect 34698 4088 34704 4140
rect 34756 4088 34762 4140
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 34885 4131 34943 4137
rect 34885 4128 34897 4131
rect 34848 4100 34897 4128
rect 34848 4088 34854 4100
rect 34885 4097 34897 4100
rect 34931 4097 34943 4131
rect 34992 4128 35020 4168
rect 43990 4156 43996 4208
rect 44048 4196 44054 4208
rect 49418 4196 49424 4208
rect 44048 4168 49424 4196
rect 44048 4156 44054 4168
rect 49418 4156 49424 4168
rect 49476 4156 49482 4208
rect 49510 4156 49516 4208
rect 49568 4196 49574 4208
rect 49568 4168 53236 4196
rect 49568 4156 49574 4168
rect 53208 4128 53236 4168
rect 53282 4156 53288 4208
rect 53340 4196 53346 4208
rect 70486 4196 70492 4208
rect 53340 4168 70492 4196
rect 53340 4156 53346 4168
rect 70486 4156 70492 4168
rect 70544 4156 70550 4208
rect 56410 4128 56416 4140
rect 34992 4100 51074 4128
rect 53208 4100 56416 4128
rect 34885 4091 34943 4097
rect 41690 4060 41696 4072
rect 29840 4032 41696 4060
rect 41690 4020 41696 4032
rect 41748 4020 41754 4072
rect 42610 4020 42616 4072
rect 42668 4060 42674 4072
rect 46934 4060 46940 4072
rect 42668 4032 46940 4060
rect 42668 4020 42674 4032
rect 46934 4020 46940 4032
rect 46992 4020 46998 4072
rect 51046 4060 51074 4100
rect 56410 4088 56416 4100
rect 56468 4088 56474 4140
rect 61102 4088 61108 4140
rect 61160 4128 61166 4140
rect 67542 4128 67548 4140
rect 61160 4100 67548 4128
rect 61160 4088 61166 4100
rect 67542 4088 67548 4100
rect 67600 4088 67606 4140
rect 64966 4060 64972 4072
rect 51046 4032 64972 4060
rect 64966 4020 64972 4032
rect 65024 4020 65030 4072
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 40402 3992 40408 4004
rect 17920 3964 40408 3992
rect 17920 3952 17926 3964
rect 40402 3952 40408 3964
rect 40460 3952 40466 4004
rect 42518 3952 42524 4004
rect 42576 3992 42582 4004
rect 45094 3992 45100 4004
rect 42576 3964 45100 3992
rect 42576 3952 42582 3964
rect 45094 3952 45100 3964
rect 45152 3952 45158 4004
rect 54018 3952 54024 4004
rect 54076 3992 54082 4004
rect 54570 3992 54576 4004
rect 54076 3964 54576 3992
rect 54076 3952 54082 3964
rect 54570 3952 54576 3964
rect 54628 3952 54634 4004
rect 60826 3952 60832 4004
rect 60884 3992 60890 4004
rect 62758 3992 62764 4004
rect 60884 3964 62764 3992
rect 60884 3952 60890 3964
rect 62758 3952 62764 3964
rect 62816 3952 62822 4004
rect 23566 3884 23572 3936
rect 23624 3924 23630 3936
rect 27614 3924 27620 3936
rect 23624 3896 27620 3924
rect 23624 3884 23630 3896
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 27706 3884 27712 3936
rect 27764 3884 27770 3936
rect 30377 3927 30435 3933
rect 30377 3893 30389 3927
rect 30423 3924 30435 3927
rect 33962 3924 33968 3936
rect 30423 3896 33968 3924
rect 30423 3893 30435 3896
rect 30377 3887 30435 3893
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 49142 3924 49148 3936
rect 36044 3896 49148 3924
rect 36044 3884 36050 3896
rect 49142 3884 49148 3896
rect 49200 3884 49206 3936
rect 1012 3834 74980 3856
rect 1012 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 74980 3834
rect 1012 3760 74980 3782
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 26050 3680 26056 3732
rect 26108 3680 26114 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 29730 3720 29736 3732
rect 26283 3692 29736 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 29730 3680 29736 3692
rect 29788 3680 29794 3732
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 31389 3723 31447 3729
rect 31389 3720 31401 3723
rect 31352 3692 31401 3720
rect 31352 3680 31358 3692
rect 31389 3689 31401 3692
rect 31435 3689 31447 3723
rect 31389 3683 31447 3689
rect 32398 3680 32404 3732
rect 32456 3680 32462 3732
rect 33152 3692 33364 3720
rect 33152 3652 33180 3692
rect 19444 3624 25268 3652
rect 19444 3593 19472 3624
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3553 19487 3587
rect 19429 3547 19487 3553
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 20680 3556 23673 3584
rect 20680 3544 20686 3556
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 24946 3544 24952 3596
rect 25004 3544 25010 3596
rect 25240 3584 25268 3624
rect 25424 3624 33180 3652
rect 33336 3652 33364 3692
rect 33410 3680 33416 3732
rect 33468 3720 33474 3732
rect 47486 3720 47492 3732
rect 33468 3692 47492 3720
rect 33468 3680 33474 3692
rect 47486 3680 47492 3692
rect 47544 3680 47550 3732
rect 58526 3680 58532 3732
rect 58584 3720 58590 3732
rect 61286 3720 61292 3732
rect 58584 3692 61292 3720
rect 58584 3680 58590 3692
rect 61286 3680 61292 3692
rect 61344 3680 61350 3732
rect 41230 3652 41236 3664
rect 33336 3624 41236 3652
rect 25424 3584 25452 3624
rect 41230 3612 41236 3624
rect 41288 3612 41294 3664
rect 42242 3612 42248 3664
rect 42300 3652 42306 3664
rect 52638 3652 52644 3664
rect 42300 3624 52644 3652
rect 42300 3612 42306 3624
rect 52638 3612 52644 3624
rect 52696 3612 52702 3664
rect 55766 3612 55772 3664
rect 55824 3652 55830 3664
rect 66254 3652 66260 3664
rect 55824 3624 66260 3652
rect 55824 3612 55830 3624
rect 66254 3612 66260 3624
rect 66312 3612 66318 3664
rect 25240 3556 25452 3584
rect 25593 3587 25651 3593
rect 25593 3553 25605 3587
rect 25639 3584 25651 3587
rect 28810 3584 28816 3596
rect 25639 3556 28816 3584
rect 25639 3553 25651 3556
rect 25593 3547 25651 3553
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 31386 3584 31392 3596
rect 31128 3556 31392 3584
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19153 3519 19211 3525
rect 19153 3516 19165 3519
rect 18288 3488 19165 3516
rect 18288 3476 18294 3488
rect 19153 3485 19165 3488
rect 19199 3485 19211 3519
rect 19153 3479 19211 3485
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20530 3516 20536 3528
rect 20211 3488 20536 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22520 3488 22569 3516
rect 22520 3476 22526 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23566 3516 23572 3528
rect 23523 3488 23572 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 25222 3476 25228 3528
rect 25280 3476 25286 3528
rect 25774 3476 25780 3528
rect 25832 3476 25838 3528
rect 27982 3516 27988 3528
rect 25976 3488 27988 3516
rect 19889 3451 19947 3457
rect 19889 3417 19901 3451
rect 19935 3448 19947 3451
rect 19935 3420 24440 3448
rect 19935 3417 19947 3420
rect 19889 3411 19947 3417
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 23201 3383 23259 3389
rect 23201 3380 23213 3383
rect 23164 3352 23213 3380
rect 23164 3340 23170 3352
rect 23201 3349 23213 3352
rect 23247 3349 23259 3383
rect 23201 3343 23259 3349
rect 23290 3340 23296 3392
rect 23348 3340 23354 3392
rect 24412 3380 24440 3420
rect 25866 3408 25872 3460
rect 25924 3408 25930 3460
rect 25976 3380 26004 3488
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 28077 3519 28135 3525
rect 28077 3485 28089 3519
rect 28123 3516 28135 3519
rect 28718 3516 28724 3528
rect 28123 3488 28724 3516
rect 28123 3485 28135 3488
rect 28077 3479 28135 3485
rect 28718 3476 28724 3488
rect 28776 3476 28782 3528
rect 31128 3516 31156 3556
rect 31386 3544 31392 3556
rect 31444 3544 31450 3596
rect 31496 3556 31892 3584
rect 28828 3488 31156 3516
rect 26142 3457 26148 3460
rect 26085 3451 26148 3457
rect 26085 3417 26097 3451
rect 26131 3417 26148 3451
rect 26085 3411 26148 3417
rect 26142 3408 26148 3411
rect 26200 3408 26206 3460
rect 27706 3408 27712 3460
rect 27764 3408 27770 3460
rect 28166 3408 28172 3460
rect 28224 3448 28230 3460
rect 28828 3448 28856 3488
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 28224 3420 28856 3448
rect 28224 3408 28230 3420
rect 28994 3408 29000 3460
rect 29052 3448 29058 3460
rect 31496 3448 31524 3556
rect 31662 3476 31668 3528
rect 31720 3476 31726 3528
rect 29052 3420 31524 3448
rect 31864 3448 31892 3556
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 39758 3584 39764 3596
rect 32456 3556 39764 3584
rect 32456 3544 32462 3556
rect 39758 3544 39764 3556
rect 39816 3544 39822 3596
rect 51534 3544 51540 3596
rect 51592 3584 51598 3596
rect 66346 3584 66352 3596
rect 51592 3556 66352 3584
rect 51592 3544 51598 3556
rect 66346 3544 66352 3556
rect 66404 3544 66410 3596
rect 32214 3476 32220 3528
rect 32272 3476 32278 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32861 3519 32919 3525
rect 32364 3512 32812 3516
rect 32861 3512 32873 3519
rect 32364 3488 32873 3512
rect 32364 3476 32370 3488
rect 32784 3485 32873 3488
rect 32907 3485 32919 3519
rect 32784 3484 32919 3485
rect 32861 3479 32919 3484
rect 33042 3476 33048 3528
rect 33100 3516 33106 3528
rect 38010 3516 38016 3528
rect 33100 3488 38016 3516
rect 33100 3476 33106 3488
rect 38010 3476 38016 3488
rect 38068 3476 38074 3528
rect 44818 3476 44824 3528
rect 44876 3516 44882 3528
rect 58526 3516 58532 3528
rect 44876 3488 58532 3516
rect 44876 3476 44882 3488
rect 58526 3476 58532 3488
rect 58584 3476 58590 3528
rect 60734 3476 60740 3528
rect 60792 3516 60798 3528
rect 67082 3516 67088 3528
rect 60792 3488 67088 3516
rect 60792 3476 60798 3488
rect 67082 3476 67088 3488
rect 67140 3476 67146 3528
rect 44634 3448 44640 3460
rect 31864 3420 44640 3448
rect 29052 3408 29058 3420
rect 44634 3408 44640 3420
rect 44692 3408 44698 3460
rect 48222 3408 48228 3460
rect 48280 3448 48286 3460
rect 66990 3448 66996 3460
rect 48280 3420 66996 3448
rect 48280 3408 48286 3420
rect 66990 3408 66996 3420
rect 67048 3408 67054 3460
rect 24412 3352 26004 3380
rect 27617 3383 27675 3389
rect 27617 3349 27629 3383
rect 27663 3380 27675 3383
rect 27798 3380 27804 3392
rect 27663 3352 27804 3380
rect 27663 3349 27675 3352
rect 27617 3343 27675 3349
rect 27798 3340 27804 3352
rect 27856 3340 27862 3392
rect 27890 3340 27896 3392
rect 27948 3340 27954 3392
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 31018 3380 31024 3392
rect 28040 3352 31024 3380
rect 28040 3340 28046 3352
rect 31018 3340 31024 3352
rect 31076 3340 31082 3392
rect 31849 3383 31907 3389
rect 31849 3349 31861 3383
rect 31895 3380 31907 3383
rect 32674 3380 32680 3392
rect 31895 3352 32680 3380
rect 31895 3349 31907 3352
rect 31849 3343 31907 3349
rect 32674 3340 32680 3352
rect 32732 3340 32738 3392
rect 33045 3383 33103 3389
rect 33045 3349 33057 3383
rect 33091 3380 33103 3383
rect 36906 3380 36912 3392
rect 33091 3352 36912 3380
rect 33091 3349 33103 3352
rect 33045 3343 33103 3349
rect 36906 3340 36912 3352
rect 36964 3340 36970 3392
rect 36998 3340 37004 3392
rect 37056 3380 37062 3392
rect 47486 3380 47492 3392
rect 37056 3352 47492 3380
rect 37056 3340 37062 3352
rect 47486 3340 47492 3352
rect 47544 3340 47550 3392
rect 1012 3290 74980 3312
rect 1012 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74980 3290
rect 1012 3216 74980 3238
rect 20530 3136 20536 3188
rect 20588 3136 20594 3188
rect 20898 3136 20904 3188
rect 20956 3136 20962 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 24854 3176 24860 3188
rect 21315 3148 24860 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 25774 3136 25780 3188
rect 25832 3176 25838 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25832 3148 25881 3176
rect 25832 3136 25838 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 27706 3136 27712 3188
rect 27764 3176 27770 3188
rect 28077 3179 28135 3185
rect 28077 3176 28089 3179
rect 27764 3148 28089 3176
rect 27764 3136 27770 3148
rect 28077 3145 28089 3148
rect 28123 3145 28135 3179
rect 28077 3139 28135 3145
rect 29457 3179 29515 3185
rect 29457 3145 29469 3179
rect 29503 3176 29515 3179
rect 29546 3176 29552 3188
rect 29503 3148 29552 3176
rect 29503 3145 29515 3148
rect 29457 3139 29515 3145
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 30193 3179 30251 3185
rect 30193 3145 30205 3179
rect 30239 3145 30251 3179
rect 30193 3139 30251 3145
rect 31481 3179 31539 3185
rect 31481 3145 31493 3179
rect 31527 3176 31539 3179
rect 33410 3176 33416 3188
rect 31527 3148 33416 3176
rect 31527 3145 31539 3148
rect 31481 3139 31539 3145
rect 17862 3068 17868 3120
rect 17920 3068 17926 3120
rect 21110 3111 21168 3117
rect 21110 3077 21122 3111
rect 21156 3108 21168 3111
rect 22830 3108 22836 3120
rect 21156 3080 22836 3108
rect 21156 3077 21168 3080
rect 21110 3071 21168 3077
rect 22830 3068 22836 3080
rect 22888 3068 22894 3120
rect 26050 3108 26056 3120
rect 22940 3080 26056 3108
rect 18138 3000 18144 3052
rect 18196 3000 18202 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 20622 3040 20628 3052
rect 19392 3012 20628 3040
rect 19392 3000 19398 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 20772 3012 21373 3040
rect 20772 3000 20778 3012
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 21468 3012 22094 3040
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 18969 2975 19027 2981
rect 18969 2972 18981 2975
rect 18748 2944 18981 2972
rect 18748 2932 18754 2944
rect 18969 2941 18981 2944
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 19150 2932 19156 2984
rect 19208 2932 19214 2984
rect 19886 2932 19892 2984
rect 19944 2932 19950 2984
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2972 21051 2975
rect 21468 2972 21496 3012
rect 21039 2944 21496 2972
rect 21039 2941 21051 2944
rect 20993 2935 21051 2941
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 21008 2904 21036 2935
rect 21726 2932 21732 2984
rect 21784 2932 21790 2984
rect 22066 2972 22094 3012
rect 22940 2972 22968 3080
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 29362 3108 29368 3120
rect 26712 3080 29368 3108
rect 23106 3000 23112 3052
rect 23164 3000 23170 3052
rect 26712 3049 26740 3080
rect 29362 3068 29368 3080
rect 29420 3068 29426 3120
rect 30208 3108 30236 3139
rect 33410 3136 33416 3148
rect 33468 3136 33474 3188
rect 33505 3179 33563 3185
rect 33505 3145 33517 3179
rect 33551 3176 33563 3179
rect 33551 3148 35664 3176
rect 33551 3145 33563 3148
rect 33505 3139 33563 3145
rect 33226 3108 33232 3120
rect 30208 3080 33232 3108
rect 33226 3068 33232 3080
rect 33284 3068 33290 3120
rect 34790 3108 34796 3120
rect 33428 3080 34796 3108
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26697 3043 26755 3049
rect 26191 3012 26648 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 22066 2944 22968 2972
rect 23014 2932 23020 2984
rect 23072 2972 23078 2984
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 23072 2944 23765 2972
rect 23072 2932 23078 2944
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 24026 2932 24032 2984
rect 24084 2972 24090 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 24084 2944 24317 2972
rect 24084 2932 24090 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 25314 2932 25320 2984
rect 25372 2932 25378 2984
rect 20680 2876 21036 2904
rect 20680 2864 20686 2876
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 22336 2876 22477 2904
rect 22336 2864 22342 2876
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22465 2867 22523 2873
rect 22830 2864 22836 2916
rect 22888 2904 22894 2916
rect 26142 2904 26148 2916
rect 22888 2876 26148 2904
rect 22888 2864 22894 2876
rect 26142 2864 26148 2876
rect 26200 2864 26206 2916
rect 26620 2904 26648 3012
rect 26697 3009 26709 3043
rect 26743 3009 26755 3043
rect 26697 3003 26755 3009
rect 26881 3043 26939 3049
rect 26881 3009 26893 3043
rect 26927 3040 26939 3043
rect 26970 3040 26976 3052
rect 26927 3012 26976 3040
rect 26927 3009 26939 3012
rect 26881 3003 26939 3009
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 28534 3000 28540 3052
rect 28592 3000 28598 3052
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 28960 3012 29040 3040
rect 28960 3000 28966 3012
rect 27062 2932 27068 2984
rect 27120 2932 27126 2984
rect 27522 2932 27528 2984
rect 27580 2932 27586 2984
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 28813 2975 28871 2981
rect 28813 2972 28825 2975
rect 28776 2944 28825 2972
rect 28776 2932 28782 2944
rect 28813 2941 28825 2944
rect 28859 2941 28871 2975
rect 29012 2972 29040 3012
rect 29086 3000 29092 3052
rect 29144 3000 29150 3052
rect 29546 3000 29552 3052
rect 29604 3000 29610 3052
rect 29638 3000 29644 3052
rect 29696 3040 29702 3052
rect 29733 3043 29791 3049
rect 29733 3040 29745 3043
rect 29696 3012 29745 3040
rect 29696 3000 29702 3012
rect 29733 3009 29745 3012
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 30006 3000 30012 3052
rect 30064 3000 30070 3052
rect 31570 3000 31576 3052
rect 31628 3000 31634 3052
rect 32033 3043 32091 3049
rect 32033 3009 32045 3043
rect 32079 3040 32091 3043
rect 32306 3040 32312 3052
rect 32079 3012 32312 3040
rect 32079 3009 32091 3012
rect 32033 3003 32091 3009
rect 32306 3000 32312 3012
rect 32364 3000 32370 3052
rect 32582 3000 32588 3052
rect 32640 3000 32646 3052
rect 32953 3043 33011 3049
rect 32953 3009 32965 3043
rect 32999 3040 33011 3043
rect 33134 3040 33140 3052
rect 32999 3012 33140 3040
rect 32999 3009 33011 3012
rect 32953 3003 33011 3009
rect 33134 3000 33140 3012
rect 33192 3000 33198 3052
rect 33318 3000 33324 3052
rect 33376 3000 33382 3052
rect 29012 2944 29592 2972
rect 28813 2935 28871 2941
rect 29454 2904 29460 2916
rect 26620 2876 29460 2904
rect 29454 2864 29460 2876
rect 29512 2864 29518 2916
rect 18414 2796 18420 2848
rect 18472 2796 18478 2848
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 21450 2796 21456 2848
rect 21508 2796 21514 2848
rect 22370 2796 22376 2848
rect 22428 2796 22434 2848
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 23201 2839 23259 2845
rect 23201 2836 23213 2839
rect 22612 2808 23213 2836
rect 22612 2796 22618 2808
rect 23201 2805 23213 2808
rect 23247 2805 23259 2839
rect 23201 2799 23259 2805
rect 24946 2796 24952 2848
rect 25004 2796 25010 2848
rect 25958 2796 25964 2848
rect 26016 2796 26022 2848
rect 26510 2796 26516 2848
rect 26568 2796 26574 2848
rect 28074 2796 28080 2848
rect 28132 2836 28138 2848
rect 28353 2839 28411 2845
rect 28353 2836 28365 2839
rect 28132 2808 28365 2836
rect 28132 2796 28138 2808
rect 28353 2805 28365 2808
rect 28399 2805 28411 2839
rect 29564 2836 29592 2944
rect 30190 2932 30196 2984
rect 30248 2972 30254 2984
rect 30285 2975 30343 2981
rect 30285 2972 30297 2975
rect 30248 2944 30297 2972
rect 30248 2932 30254 2944
rect 30285 2941 30297 2944
rect 30331 2941 30343 2975
rect 30285 2935 30343 2941
rect 30926 2932 30932 2984
rect 30984 2932 30990 2984
rect 32214 2932 32220 2984
rect 32272 2932 32278 2984
rect 33428 2972 33456 3080
rect 34790 3068 34796 3080
rect 34848 3068 34854 3120
rect 33778 3000 33784 3052
rect 33836 3000 33842 3052
rect 34054 3000 34060 3052
rect 34112 3000 34118 3052
rect 34517 3043 34575 3049
rect 34517 3009 34529 3043
rect 34563 3040 34575 3043
rect 34606 3040 34612 3052
rect 34563 3012 34612 3040
rect 34563 3009 34575 3012
rect 34517 3003 34575 3009
rect 34606 3000 34612 3012
rect 34664 3000 34670 3052
rect 34882 3000 34888 3052
rect 34940 3000 34946 3052
rect 35161 2975 35219 2981
rect 35161 2972 35173 2975
rect 32508 2944 33456 2972
rect 33980 2944 35173 2972
rect 29917 2907 29975 2913
rect 29917 2873 29929 2907
rect 29963 2904 29975 2907
rect 32508 2904 32536 2944
rect 33980 2904 34008 2944
rect 35161 2941 35173 2944
rect 35207 2941 35219 2975
rect 35636 2972 35664 3148
rect 36998 3136 37004 3188
rect 37056 3136 37062 3188
rect 35897 3111 35955 3117
rect 35897 3077 35909 3111
rect 35943 3108 35955 3111
rect 35986 3108 35992 3120
rect 35943 3080 35992 3108
rect 35943 3077 35955 3080
rect 35897 3071 35955 3077
rect 35986 3068 35992 3080
rect 36044 3068 36050 3120
rect 47026 3068 47032 3120
rect 47084 3108 47090 3120
rect 51258 3108 51264 3120
rect 47084 3080 51264 3108
rect 47084 3068 47090 3080
rect 51258 3068 51264 3080
rect 51316 3068 51322 3120
rect 54573 3111 54631 3117
rect 54573 3077 54585 3111
rect 54619 3108 54631 3111
rect 63954 3108 63960 3120
rect 54619 3080 63960 3108
rect 54619 3077 54631 3080
rect 54573 3071 54631 3077
rect 63954 3068 63960 3080
rect 64012 3068 64018 3120
rect 35710 3000 35716 3052
rect 35768 3000 35774 3052
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 36722 3040 36728 3052
rect 36311 3012 36728 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 36722 3000 36728 3012
rect 36780 3000 36786 3052
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 36906 3000 36912 3052
rect 36964 3040 36970 3052
rect 42426 3040 42432 3052
rect 36964 3012 42432 3040
rect 36964 3000 36970 3012
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45922 3000 45928 3052
rect 45980 3000 45986 3052
rect 47118 3000 47124 3052
rect 47176 3040 47182 3052
rect 47489 3043 47547 3049
rect 47489 3040 47501 3043
rect 47176 3012 47501 3040
rect 47176 3000 47182 3012
rect 47489 3009 47501 3012
rect 47535 3009 47547 3043
rect 47489 3003 47547 3009
rect 49050 3000 49056 3052
rect 49108 3000 49114 3052
rect 52914 3000 52920 3052
rect 52972 3000 52978 3052
rect 53926 3000 53932 3052
rect 53984 3040 53990 3052
rect 54205 3043 54263 3049
rect 54205 3040 54217 3043
rect 53984 3012 54217 3040
rect 53984 3000 53990 3012
rect 54205 3009 54217 3012
rect 54251 3009 54263 3043
rect 54205 3003 54263 3009
rect 54662 3000 54668 3052
rect 54720 3000 54726 3052
rect 56226 3000 56232 3052
rect 56284 3000 56290 3052
rect 57790 3000 57796 3052
rect 57848 3000 57854 3052
rect 59446 3000 59452 3052
rect 59504 3000 59510 3052
rect 61194 3000 61200 3052
rect 61252 3000 61258 3052
rect 63218 3000 63224 3052
rect 63276 3000 63282 3052
rect 64782 3000 64788 3052
rect 64840 3000 64846 3052
rect 66438 3000 66444 3052
rect 66496 3000 66502 3052
rect 68094 3000 68100 3052
rect 68152 3000 68158 3052
rect 69842 3000 69848 3052
rect 69900 3000 69906 3052
rect 71406 3000 71412 3052
rect 71464 3000 71470 3052
rect 72881 3043 72939 3049
rect 72881 3009 72893 3043
rect 72927 3040 72939 3043
rect 73246 3040 73252 3052
rect 72927 3012 73252 3040
rect 72927 3009 72939 3012
rect 72881 3003 72939 3009
rect 73246 3000 73252 3012
rect 73304 3000 73310 3052
rect 42978 2972 42984 2984
rect 35636 2944 42984 2972
rect 35161 2935 35219 2941
rect 42978 2932 42984 2944
rect 43036 2932 43042 2984
rect 29963 2876 32536 2904
rect 32600 2876 34008 2904
rect 35069 2907 35127 2913
rect 29963 2873 29975 2876
rect 29917 2867 29975 2873
rect 32600 2836 32628 2876
rect 35069 2873 35081 2907
rect 35115 2873 35127 2907
rect 35069 2867 35127 2873
rect 29564 2808 32628 2836
rect 28353 2799 28411 2805
rect 33870 2796 33876 2848
rect 33928 2836 33934 2848
rect 34241 2839 34299 2845
rect 34241 2836 34253 2839
rect 33928 2808 34253 2836
rect 33928 2796 33934 2808
rect 34241 2805 34253 2808
rect 34287 2805 34299 2839
rect 35084 2836 35112 2867
rect 35710 2864 35716 2916
rect 35768 2904 35774 2916
rect 44818 2904 44824 2916
rect 35768 2876 44824 2904
rect 35768 2864 35774 2876
rect 44818 2864 44824 2876
rect 44876 2864 44882 2916
rect 47673 2907 47731 2913
rect 47673 2873 47685 2907
rect 47719 2904 47731 2907
rect 50062 2904 50068 2916
rect 47719 2876 50068 2904
rect 47719 2873 47731 2876
rect 47673 2867 47731 2873
rect 50062 2864 50068 2876
rect 50120 2864 50126 2916
rect 44910 2836 44916 2848
rect 35084 2808 44916 2836
rect 34241 2799 34299 2805
rect 44910 2796 44916 2808
rect 44968 2796 44974 2848
rect 46109 2839 46167 2845
rect 46109 2805 46121 2839
rect 46155 2836 46167 2839
rect 47578 2836 47584 2848
rect 46155 2808 47584 2836
rect 46155 2805 46167 2808
rect 46109 2799 46167 2805
rect 47578 2796 47584 2808
rect 47636 2796 47642 2848
rect 49237 2839 49295 2845
rect 49237 2805 49249 2839
rect 49283 2836 49295 2839
rect 52638 2836 52644 2848
rect 49283 2808 52644 2836
rect 49283 2805 49295 2808
rect 49237 2799 49295 2805
rect 52638 2796 52644 2808
rect 52696 2796 52702 2848
rect 53098 2796 53104 2848
rect 53156 2796 53162 2848
rect 54849 2839 54907 2845
rect 54849 2805 54861 2839
rect 54895 2836 54907 2839
rect 55214 2836 55220 2848
rect 54895 2808 55220 2836
rect 54895 2805 54907 2808
rect 54849 2799 54907 2805
rect 55214 2796 55220 2808
rect 55272 2796 55278 2848
rect 56410 2796 56416 2848
rect 56468 2796 56474 2848
rect 57974 2796 57980 2848
rect 58032 2796 58038 2848
rect 59633 2839 59691 2845
rect 59633 2805 59645 2839
rect 59679 2836 59691 2839
rect 60366 2836 60372 2848
rect 59679 2808 60372 2836
rect 59679 2805 59691 2808
rect 59633 2799 59691 2805
rect 60366 2796 60372 2808
rect 60424 2796 60430 2848
rect 61378 2796 61384 2848
rect 61436 2796 61442 2848
rect 63034 2796 63040 2848
rect 63092 2796 63098 2848
rect 64598 2796 64604 2848
rect 64656 2796 64662 2848
rect 66254 2796 66260 2848
rect 66312 2796 66318 2848
rect 68278 2796 68284 2848
rect 68336 2796 68342 2848
rect 69658 2796 69664 2848
rect 69716 2796 69722 2848
rect 71222 2796 71228 2848
rect 71280 2796 71286 2848
rect 73065 2839 73123 2845
rect 73065 2805 73077 2839
rect 73111 2836 73123 2839
rect 73246 2836 73252 2848
rect 73111 2808 73252 2836
rect 73111 2805 73123 2808
rect 73065 2799 73123 2805
rect 73246 2796 73252 2808
rect 73304 2796 73310 2848
rect 1012 2746 74980 2768
rect 1012 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 74980 2746
rect 1012 2672 74980 2694
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 18196 2604 18245 2632
rect 18196 2592 18202 2604
rect 18233 2601 18245 2604
rect 18279 2601 18291 2635
rect 18233 2595 18291 2601
rect 18969 2635 19027 2641
rect 18969 2601 18981 2635
rect 19015 2632 19027 2635
rect 19150 2632 19156 2644
rect 19015 2604 19156 2632
rect 19015 2601 19027 2604
rect 18969 2595 19027 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19886 2592 19892 2644
rect 19944 2592 19950 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20806 2632 20812 2644
rect 20027 2604 20812 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 21361 2635 21419 2641
rect 21361 2601 21373 2635
rect 21407 2632 21419 2635
rect 21726 2632 21732 2644
rect 21407 2604 21732 2632
rect 21407 2601 21419 2604
rect 21361 2595 21419 2601
rect 21726 2592 21732 2604
rect 21784 2592 21790 2644
rect 23290 2632 23296 2644
rect 21836 2604 23296 2632
rect 21836 2564 21864 2604
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 24026 2592 24032 2644
rect 24084 2632 24090 2644
rect 24121 2635 24179 2641
rect 24121 2632 24133 2635
rect 24084 2604 24133 2632
rect 24084 2592 24090 2604
rect 24121 2601 24133 2604
rect 24167 2601 24179 2635
rect 24121 2595 24179 2601
rect 25222 2592 25228 2644
rect 25280 2592 25286 2644
rect 25314 2592 25320 2644
rect 25372 2592 25378 2644
rect 27522 2592 27528 2644
rect 27580 2592 27586 2644
rect 29086 2592 29092 2644
rect 29144 2632 29150 2644
rect 29273 2635 29331 2641
rect 29273 2632 29285 2635
rect 29144 2604 29285 2632
rect 29144 2592 29150 2604
rect 29273 2601 29285 2604
rect 29319 2601 29331 2635
rect 29273 2595 29331 2601
rect 31570 2592 31576 2644
rect 31628 2632 31634 2644
rect 31665 2635 31723 2641
rect 31665 2632 31677 2635
rect 31628 2604 31677 2632
rect 31628 2592 31634 2604
rect 31665 2601 31677 2604
rect 31711 2601 31723 2635
rect 31665 2595 31723 2601
rect 33134 2592 33140 2644
rect 33192 2592 33198 2644
rect 34054 2592 34060 2644
rect 34112 2632 34118 2644
rect 34241 2635 34299 2641
rect 34241 2632 34253 2635
rect 34112 2604 34253 2632
rect 34112 2592 34118 2604
rect 34241 2601 34253 2604
rect 34287 2601 34299 2635
rect 34241 2595 34299 2601
rect 36170 2592 36176 2644
rect 36228 2632 36234 2644
rect 46566 2632 46572 2644
rect 36228 2604 46572 2632
rect 36228 2592 36234 2604
rect 46566 2592 46572 2604
rect 46624 2592 46630 2644
rect 47121 2635 47179 2641
rect 47121 2601 47133 2635
rect 47167 2632 47179 2635
rect 48222 2632 48228 2644
rect 47167 2604 48228 2632
rect 47167 2601 47179 2604
rect 47121 2595 47179 2601
rect 48222 2592 48228 2604
rect 48280 2592 48286 2644
rect 53926 2592 53932 2644
rect 53984 2592 53990 2644
rect 56045 2635 56103 2641
rect 56045 2601 56057 2635
rect 56091 2632 56103 2635
rect 60734 2632 60740 2644
rect 56091 2604 60740 2632
rect 56091 2601 56103 2604
rect 56045 2595 56103 2601
rect 60734 2592 60740 2604
rect 60792 2592 60798 2644
rect 63313 2635 63371 2641
rect 63313 2601 63325 2635
rect 63359 2632 63371 2635
rect 67358 2632 67364 2644
rect 63359 2604 67364 2632
rect 63359 2601 63371 2604
rect 63313 2595 63371 2601
rect 67358 2592 67364 2604
rect 67416 2592 67422 2644
rect 17512 2536 21864 2564
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17512 2437 17540 2536
rect 25866 2524 25872 2576
rect 25924 2564 25930 2576
rect 30466 2564 30472 2576
rect 25924 2536 30472 2564
rect 25924 2524 25930 2536
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 30576 2536 35894 2564
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2496 18475 2499
rect 19702 2496 19708 2508
rect 18463 2468 19708 2496
rect 18463 2465 18475 2468
rect 18417 2459 18475 2465
rect 19702 2456 19708 2468
rect 19760 2456 19766 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 20806 2496 20812 2508
rect 20671 2468 20812 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 25958 2496 25964 2508
rect 22848 2468 25964 2496
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 17000 2400 17049 2428
rect 17000 2388 17006 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 19337 2431 19395 2437
rect 19337 2397 19349 2431
rect 19383 2428 19395 2431
rect 20254 2428 20260 2440
rect 19383 2400 20260 2428
rect 19383 2397 19395 2400
rect 19337 2391 19395 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20622 2360 20628 2372
rect 17236 2332 20628 2360
rect 17236 2301 17264 2332
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 20732 2360 20760 2391
rect 21358 2388 21364 2440
rect 21416 2428 21422 2440
rect 22848 2437 22876 2468
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 28442 2456 28448 2508
rect 28500 2496 28506 2508
rect 30576 2496 30604 2536
rect 28500 2468 30604 2496
rect 28500 2456 28506 2468
rect 30926 2456 30932 2508
rect 30984 2456 30990 2508
rect 35866 2496 35894 2536
rect 39298 2524 39304 2576
rect 39356 2524 39362 2576
rect 44361 2567 44419 2573
rect 44361 2533 44373 2567
rect 44407 2564 44419 2567
rect 44726 2564 44732 2576
rect 44407 2536 44732 2564
rect 44407 2533 44419 2536
rect 44361 2527 44419 2533
rect 44726 2524 44732 2536
rect 44784 2524 44790 2576
rect 47210 2524 47216 2576
rect 47268 2564 47274 2576
rect 55306 2564 55312 2576
rect 47268 2536 55312 2564
rect 47268 2524 47274 2536
rect 55306 2524 55312 2536
rect 55364 2524 55370 2576
rect 68738 2564 68744 2576
rect 60016 2536 68744 2564
rect 60016 2496 60044 2536
rect 68738 2524 68744 2536
rect 68796 2524 68802 2576
rect 35866 2468 60044 2496
rect 60737 2499 60795 2505
rect 60737 2465 60749 2499
rect 60783 2496 60795 2499
rect 65794 2496 65800 2508
rect 60783 2468 65800 2496
rect 60783 2465 60795 2468
rect 60737 2459 60795 2465
rect 65794 2456 65800 2468
rect 65852 2456 65858 2508
rect 67450 2456 67456 2508
rect 67508 2456 67514 2508
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 21416 2400 21649 2428
rect 21416 2388 21422 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 24026 2428 24032 2440
rect 23615 2400 24032 2428
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25280 2400 25881 2428
rect 25280 2388 25286 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26050 2388 26056 2440
rect 26108 2388 26114 2440
rect 26878 2388 26884 2440
rect 26936 2428 26942 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26936 2400 27353 2428
rect 26936 2388 26942 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27430 2388 27436 2440
rect 27488 2428 27494 2440
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 27488 2400 28089 2428
rect 27488 2388 27494 2400
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28258 2388 28264 2440
rect 28316 2428 28322 2440
rect 28353 2431 28411 2437
rect 28353 2428 28365 2431
rect 28316 2400 28365 2428
rect 28316 2388 28322 2400
rect 28353 2397 28365 2400
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28626 2388 28632 2440
rect 28684 2388 28690 2440
rect 29178 2388 29184 2440
rect 29236 2428 29242 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29236 2400 30021 2428
rect 29236 2388 29242 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 30009 2391 30067 2397
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32490 2388 32496 2440
rect 32548 2388 32554 2440
rect 33594 2388 33600 2440
rect 33652 2388 33658 2440
rect 35161 2431 35219 2437
rect 35161 2397 35173 2431
rect 35207 2428 35219 2431
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35207 2400 35265 2428
rect 35207 2397 35219 2400
rect 35161 2391 35219 2397
rect 35253 2397 35265 2400
rect 35299 2397 35311 2431
rect 35253 2391 35311 2397
rect 35897 2431 35955 2437
rect 35897 2397 35909 2431
rect 35943 2428 35955 2431
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35943 2400 36001 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36538 2388 36544 2440
rect 36596 2388 36602 2440
rect 41414 2428 41420 2440
rect 39040 2400 41420 2428
rect 21726 2360 21732 2372
rect 20732 2332 21732 2360
rect 21726 2320 21732 2332
rect 21784 2320 21790 2372
rect 23201 2363 23259 2369
rect 23201 2329 23213 2363
rect 23247 2360 23259 2363
rect 34885 2363 34943 2369
rect 23247 2332 31892 2360
rect 23247 2329 23259 2332
rect 23201 2323 23259 2329
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17313 2295 17371 2301
rect 17313 2261 17325 2295
rect 17359 2292 17371 2295
rect 17770 2292 17776 2304
rect 17359 2264 17776 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 20898 2292 20904 2304
rect 18380 2264 20904 2292
rect 18380 2252 18386 2264
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 26694 2252 26700 2304
rect 26752 2252 26758 2304
rect 26786 2252 26792 2304
rect 26844 2252 26850 2304
rect 28534 2252 28540 2304
rect 28592 2252 28598 2304
rect 29086 2252 29092 2304
rect 29144 2292 29150 2304
rect 29457 2295 29515 2301
rect 29457 2292 29469 2295
rect 29144 2264 29469 2292
rect 29144 2252 29150 2264
rect 29457 2261 29469 2264
rect 29503 2261 29515 2295
rect 29457 2255 29515 2261
rect 30282 2252 30288 2304
rect 30340 2252 30346 2304
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 31757 2295 31815 2301
rect 31757 2292 31769 2295
rect 31352 2264 31769 2292
rect 31352 2252 31358 2264
rect 31757 2261 31769 2264
rect 31803 2261 31815 2295
rect 31864 2292 31892 2332
rect 34885 2329 34897 2363
rect 34931 2360 34943 2363
rect 39040 2360 39068 2400
rect 41414 2388 41420 2400
rect 41472 2388 41478 2440
rect 42334 2388 42340 2440
rect 42392 2428 42398 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 42392 2400 42441 2428
rect 42392 2388 42398 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 43496 2400 43729 2428
rect 43496 2388 43502 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 43717 2391 43775 2397
rect 44729 2431 44787 2437
rect 44729 2397 44741 2431
rect 44775 2428 44787 2431
rect 44913 2431 44971 2437
rect 44913 2428 44925 2431
rect 44775 2400 44925 2428
rect 44775 2397 44787 2400
rect 44729 2391 44787 2397
rect 44913 2397 44925 2400
rect 44959 2397 44971 2431
rect 44913 2391 44971 2397
rect 45554 2388 45560 2440
rect 45612 2388 45618 2440
rect 46198 2388 46204 2440
rect 46256 2388 46262 2440
rect 47302 2388 47308 2440
rect 47360 2428 47366 2440
rect 47397 2431 47455 2437
rect 47397 2428 47409 2431
rect 47360 2400 47409 2428
rect 47360 2388 47366 2400
rect 47397 2397 47409 2400
rect 47443 2397 47455 2431
rect 48866 2428 48872 2440
rect 47397 2391 47455 2397
rect 47688 2400 48872 2428
rect 34931 2332 39068 2360
rect 34931 2329 34943 2332
rect 34885 2323 34943 2329
rect 39114 2320 39120 2372
rect 39172 2360 39178 2372
rect 39485 2363 39543 2369
rect 39485 2360 39497 2363
rect 39172 2332 39497 2360
rect 39172 2320 39178 2332
rect 39485 2329 39497 2332
rect 39531 2329 39543 2363
rect 39485 2323 39543 2329
rect 43073 2363 43131 2369
rect 43073 2329 43085 2363
rect 43119 2360 43131 2363
rect 44634 2360 44640 2372
rect 43119 2332 44640 2360
rect 43119 2329 43131 2332
rect 43073 2323 43131 2329
rect 44634 2320 44640 2332
rect 44692 2320 44698 2372
rect 47213 2363 47271 2369
rect 46676 2332 47164 2360
rect 43530 2292 43536 2304
rect 31864 2264 43536 2292
rect 31757 2255 31815 2261
rect 43530 2252 43536 2264
rect 43588 2252 43594 2304
rect 44545 2295 44603 2301
rect 44545 2261 44557 2295
rect 44591 2292 44603 2295
rect 46676 2292 46704 2332
rect 44591 2264 46704 2292
rect 46753 2295 46811 2301
rect 44591 2261 44603 2264
rect 44545 2255 44603 2261
rect 46753 2261 46765 2295
rect 46799 2292 46811 2295
rect 46842 2292 46848 2304
rect 46799 2264 46848 2292
rect 46799 2261 46811 2264
rect 46753 2255 46811 2261
rect 46842 2252 46848 2264
rect 46900 2252 46906 2304
rect 47136 2292 47164 2332
rect 47213 2329 47225 2363
rect 47259 2360 47271 2363
rect 47688 2360 47716 2400
rect 48866 2388 48872 2400
rect 48924 2388 48930 2440
rect 48958 2388 48964 2440
rect 49016 2428 49022 2440
rect 49053 2431 49111 2437
rect 49053 2428 49065 2431
rect 49016 2400 49065 2428
rect 49016 2388 49022 2400
rect 49053 2397 49065 2400
rect 49099 2397 49111 2431
rect 49053 2391 49111 2397
rect 53377 2431 53435 2437
rect 53377 2397 53389 2431
rect 53423 2428 53435 2431
rect 53834 2428 53840 2440
rect 53423 2400 53840 2428
rect 53423 2397 53435 2400
rect 53377 2391 53435 2397
rect 53834 2388 53840 2400
rect 53892 2388 53898 2440
rect 53926 2388 53932 2440
rect 53984 2428 53990 2440
rect 54113 2431 54171 2437
rect 54113 2428 54125 2431
rect 53984 2400 54125 2428
rect 53984 2388 53990 2400
rect 54113 2397 54125 2400
rect 54159 2397 54171 2431
rect 54113 2391 54171 2397
rect 55677 2431 55735 2437
rect 55677 2397 55689 2431
rect 55723 2428 55735 2431
rect 55723 2400 57284 2428
rect 55723 2397 55735 2400
rect 55677 2391 55735 2397
rect 54018 2360 54024 2372
rect 47259 2332 47716 2360
rect 47780 2332 54024 2360
rect 47259 2329 47271 2332
rect 47213 2323 47271 2329
rect 47780 2292 47808 2332
rect 54018 2320 54024 2332
rect 54076 2320 54082 2372
rect 55030 2320 55036 2372
rect 55088 2360 55094 2372
rect 55309 2363 55367 2369
rect 55309 2360 55321 2363
rect 55088 2332 55321 2360
rect 55088 2320 55094 2332
rect 55309 2329 55321 2332
rect 55355 2329 55367 2363
rect 55309 2323 55367 2329
rect 56137 2363 56195 2369
rect 56137 2329 56149 2363
rect 56183 2360 56195 2363
rect 56686 2360 56692 2372
rect 56183 2332 56692 2360
rect 56183 2329 56195 2332
rect 56137 2323 56195 2329
rect 56686 2320 56692 2332
rect 56744 2320 56750 2372
rect 57256 2360 57284 2400
rect 57330 2388 57336 2440
rect 57388 2388 57394 2440
rect 62298 2388 62304 2440
rect 62356 2388 62362 2440
rect 65518 2388 65524 2440
rect 65576 2428 65582 2440
rect 65613 2431 65671 2437
rect 65613 2428 65625 2431
rect 65576 2400 65625 2428
rect 65576 2388 65582 2400
rect 65613 2397 65625 2400
rect 65659 2397 65671 2431
rect 65613 2391 65671 2397
rect 67266 2388 67272 2440
rect 67324 2428 67330 2440
rect 67729 2431 67787 2437
rect 67729 2428 67741 2431
rect 67324 2400 67741 2428
rect 67324 2388 67330 2400
rect 67729 2397 67741 2400
rect 67775 2397 67787 2431
rect 67729 2391 67787 2397
rect 69934 2388 69940 2440
rect 69992 2388 69998 2440
rect 70486 2388 70492 2440
rect 70544 2428 70550 2440
rect 70673 2431 70731 2437
rect 70673 2428 70685 2431
rect 70544 2400 70685 2428
rect 70544 2388 70550 2400
rect 70673 2397 70685 2400
rect 70719 2397 70731 2431
rect 70673 2391 70731 2397
rect 57256 2332 60872 2360
rect 47136 2264 47808 2292
rect 48041 2295 48099 2301
rect 48041 2261 48053 2295
rect 48087 2292 48099 2295
rect 49418 2292 49424 2304
rect 48087 2264 49424 2292
rect 48087 2261 48099 2264
rect 48041 2255 48099 2261
rect 49418 2252 49424 2264
rect 49476 2252 49482 2304
rect 49510 2252 49516 2304
rect 49568 2292 49574 2304
rect 49697 2295 49755 2301
rect 49697 2292 49709 2295
rect 49568 2264 49709 2292
rect 49568 2252 49574 2264
rect 49697 2261 49709 2264
rect 49743 2261 49755 2295
rect 49697 2255 49755 2261
rect 54754 2252 54760 2304
rect 54812 2252 54818 2304
rect 57882 2252 57888 2304
rect 57940 2292 57946 2304
rect 57977 2295 58035 2301
rect 57977 2292 57989 2295
rect 57940 2264 57989 2292
rect 57940 2252 57946 2264
rect 57977 2261 57989 2264
rect 58023 2261 58035 2295
rect 60844 2292 60872 2332
rect 61010 2320 61016 2372
rect 61068 2320 61074 2372
rect 63405 2363 63463 2369
rect 62868 2332 63080 2360
rect 62868 2292 62896 2332
rect 60844 2264 62896 2292
rect 57977 2255 58035 2261
rect 62942 2252 62948 2304
rect 63000 2252 63006 2304
rect 63052 2292 63080 2332
rect 63405 2329 63417 2363
rect 63451 2360 63463 2363
rect 63586 2360 63592 2372
rect 63451 2332 63592 2360
rect 63451 2329 63463 2332
rect 63405 2323 63463 2329
rect 63586 2320 63592 2332
rect 63644 2320 63650 2372
rect 65150 2292 65156 2304
rect 63052 2264 65156 2292
rect 65150 2252 65156 2264
rect 65208 2252 65214 2304
rect 66070 2252 66076 2304
rect 66128 2292 66134 2304
rect 66257 2295 66315 2301
rect 66257 2292 66269 2295
rect 66128 2264 66269 2292
rect 66128 2252 66134 2264
rect 66257 2261 66269 2264
rect 66303 2261 66315 2295
rect 66257 2255 66315 2261
rect 69293 2295 69351 2301
rect 69293 2261 69305 2295
rect 69339 2292 69351 2295
rect 69382 2292 69388 2304
rect 69339 2264 69388 2292
rect 69339 2261 69351 2264
rect 69293 2255 69351 2261
rect 69382 2252 69388 2264
rect 69440 2252 69446 2304
rect 71038 2252 71044 2304
rect 71096 2292 71102 2304
rect 71317 2295 71375 2301
rect 71317 2292 71329 2295
rect 71096 2264 71329 2292
rect 71096 2252 71102 2264
rect 71317 2261 71329 2264
rect 71363 2261 71375 2295
rect 71317 2255 71375 2261
rect 1012 2202 74980 2224
rect 1012 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74980 2202
rect 1012 2128 74980 2150
rect 16393 2091 16451 2097
rect 16393 2057 16405 2091
rect 16439 2088 16451 2091
rect 17405 2091 17463 2097
rect 16439 2060 16574 2088
rect 16439 2057 16451 2060
rect 16393 2051 16451 2057
rect 16546 2020 16574 2060
rect 17405 2057 17417 2091
rect 17451 2088 17463 2091
rect 17586 2088 17592 2100
rect 17451 2060 17592 2088
rect 17451 2057 17463 2060
rect 17405 2051 17463 2057
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 18141 2091 18199 2097
rect 18141 2057 18153 2091
rect 18187 2088 18199 2091
rect 18230 2088 18236 2100
rect 18187 2060 18236 2088
rect 18187 2057 18199 2060
rect 18141 2051 18199 2057
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 21450 2088 21456 2100
rect 19352 2060 21456 2088
rect 18322 2020 18328 2032
rect 16546 1992 18328 2020
rect 18322 1980 18328 1992
rect 18380 1980 18386 2032
rect 19352 2020 19380 2060
rect 21450 2048 21456 2060
rect 21508 2048 21514 2100
rect 24121 2091 24179 2097
rect 24121 2057 24133 2091
rect 24167 2088 24179 2091
rect 24578 2088 24584 2100
rect 24167 2060 24584 2088
rect 24167 2057 24179 2060
rect 24121 2051 24179 2057
rect 24578 2048 24584 2060
rect 24636 2048 24642 2100
rect 25685 2091 25743 2097
rect 25685 2057 25697 2091
rect 25731 2057 25743 2091
rect 25685 2051 25743 2057
rect 26697 2091 26755 2097
rect 26697 2057 26709 2091
rect 26743 2088 26755 2091
rect 26970 2088 26976 2100
rect 26743 2060 26976 2088
rect 26743 2057 26755 2060
rect 26697 2051 26755 2057
rect 19274 1992 19380 2020
rect 19426 1980 19432 2032
rect 19484 2020 19490 2032
rect 20257 2023 20315 2029
rect 20257 2020 20269 2023
rect 19484 1992 20269 2020
rect 19484 1980 19490 1992
rect 20257 1989 20269 1992
rect 20303 1989 20315 2023
rect 25700 2020 25728 2051
rect 26970 2048 26976 2060
rect 27028 2048 27034 2100
rect 31849 2091 31907 2097
rect 28092 2060 31754 2088
rect 26786 2020 26792 2032
rect 20257 1983 20315 1989
rect 21468 1992 25728 2020
rect 26160 1992 26792 2020
rect 16209 1955 16267 1961
rect 16209 1921 16221 1955
rect 16255 1952 16267 1955
rect 16390 1952 16396 1964
rect 16255 1924 16396 1952
rect 16255 1921 16267 1924
rect 16209 1915 16267 1921
rect 16390 1912 16396 1924
rect 16448 1912 16454 1964
rect 17589 1955 17647 1961
rect 17589 1921 17601 1955
rect 17635 1952 17647 1955
rect 18414 1952 18420 1964
rect 17635 1924 18420 1952
rect 17635 1921 17647 1924
rect 17589 1915 17647 1921
rect 18414 1912 18420 1924
rect 18472 1912 18478 1964
rect 21468 1961 21496 1992
rect 21453 1955 21511 1961
rect 21453 1921 21465 1955
rect 21499 1921 21511 1955
rect 21453 1915 21511 1921
rect 22189 1955 22247 1961
rect 22189 1921 22201 1955
rect 22235 1952 22247 1955
rect 22370 1952 22376 1964
rect 22235 1924 22376 1952
rect 22235 1921 22247 1924
rect 22189 1915 22247 1921
rect 22370 1912 22376 1924
rect 22428 1912 22434 1964
rect 24397 1955 24455 1961
rect 24397 1921 24409 1955
rect 24443 1952 24455 1955
rect 24946 1952 24952 1964
rect 24443 1924 24952 1952
rect 24443 1921 24455 1924
rect 24397 1915 24455 1921
rect 24946 1912 24952 1924
rect 25004 1912 25010 1964
rect 25866 1912 25872 1964
rect 25924 1912 25930 1964
rect 26160 1961 26188 1992
rect 26786 1980 26792 1992
rect 26844 1980 26850 2032
rect 28092 2029 28120 2060
rect 28077 2023 28135 2029
rect 28077 1989 28089 2023
rect 28123 1989 28135 2023
rect 28077 1983 28135 1989
rect 28534 1980 28540 2032
rect 28592 2020 28598 2032
rect 31726 2020 31754 2060
rect 31849 2057 31861 2091
rect 31895 2088 31907 2091
rect 32306 2088 32312 2100
rect 31895 2060 32312 2088
rect 31895 2057 31907 2060
rect 31849 2051 31907 2057
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 32490 2048 32496 2100
rect 32548 2048 32554 2100
rect 34606 2048 34612 2100
rect 34664 2048 34670 2100
rect 34698 2048 34704 2100
rect 34756 2088 34762 2100
rect 36170 2088 36176 2100
rect 34756 2060 36176 2088
rect 34756 2048 34762 2060
rect 36170 2048 36176 2060
rect 36228 2048 36234 2100
rect 36722 2048 36728 2100
rect 36780 2088 36786 2100
rect 36817 2091 36875 2097
rect 36817 2088 36829 2091
rect 36780 2060 36829 2088
rect 36780 2048 36786 2060
rect 36817 2057 36829 2060
rect 36863 2057 36875 2091
rect 36817 2051 36875 2057
rect 39114 2048 39120 2100
rect 39172 2048 39178 2100
rect 39298 2048 39304 2100
rect 39356 2088 39362 2100
rect 41690 2088 41696 2100
rect 39356 2060 41696 2088
rect 39356 2048 39362 2060
rect 41690 2048 41696 2060
rect 41748 2048 41754 2100
rect 41969 2091 42027 2097
rect 41969 2057 41981 2091
rect 42015 2088 42027 2091
rect 42242 2088 42248 2100
rect 42015 2060 42248 2088
rect 42015 2057 42027 2060
rect 41969 2051 42027 2057
rect 42242 2048 42248 2060
rect 42300 2048 42306 2100
rect 44729 2091 44787 2097
rect 44729 2057 44741 2091
rect 44775 2088 44787 2091
rect 44818 2088 44824 2100
rect 44775 2060 44824 2088
rect 44775 2057 44787 2060
rect 44729 2051 44787 2057
rect 44818 2048 44824 2060
rect 44876 2048 44882 2100
rect 45462 2048 45468 2100
rect 45520 2088 45526 2100
rect 50430 2088 50436 2100
rect 45520 2060 50436 2088
rect 45520 2048 45526 2060
rect 50430 2048 50436 2060
rect 50488 2048 50494 2100
rect 50525 2091 50583 2097
rect 50525 2057 50537 2091
rect 50571 2088 50583 2091
rect 51534 2088 51540 2100
rect 50571 2060 51540 2088
rect 50571 2057 50583 2060
rect 50525 2051 50583 2057
rect 51534 2048 51540 2060
rect 51592 2048 51598 2100
rect 55030 2048 55036 2100
rect 55088 2048 55094 2100
rect 58897 2091 58955 2097
rect 58897 2057 58909 2091
rect 58943 2088 58955 2091
rect 61102 2088 61108 2100
rect 58943 2060 61108 2088
rect 58943 2057 58955 2060
rect 58897 2051 58955 2057
rect 61102 2048 61108 2060
rect 61160 2048 61166 2100
rect 63586 2048 63592 2100
rect 63644 2048 63650 2100
rect 64846 2060 67128 2088
rect 64846 2020 64874 2060
rect 28592 1992 29776 2020
rect 31726 1992 64874 2020
rect 28592 1980 28598 1992
rect 26145 1955 26203 1961
rect 26145 1921 26157 1955
rect 26191 1921 26203 1955
rect 26145 1915 26203 1921
rect 26694 1912 26700 1964
rect 26752 1952 26758 1964
rect 26881 1955 26939 1961
rect 26881 1952 26893 1955
rect 26752 1924 26893 1952
rect 26752 1912 26758 1924
rect 26881 1921 26893 1924
rect 26927 1921 26939 1955
rect 26881 1915 26939 1921
rect 28905 1955 28963 1961
rect 28905 1921 28917 1955
rect 28951 1921 28963 1955
rect 28905 1915 28963 1921
rect 16853 1887 16911 1893
rect 16853 1853 16865 1887
rect 16899 1884 16911 1887
rect 18046 1884 18052 1896
rect 16899 1856 18052 1884
rect 16899 1853 16911 1856
rect 16853 1847 16911 1853
rect 18046 1844 18052 1856
rect 18104 1844 18110 1896
rect 18233 1887 18291 1893
rect 18233 1853 18245 1887
rect 18279 1884 18291 1887
rect 19334 1884 19340 1896
rect 18279 1856 19340 1884
rect 18279 1853 18291 1856
rect 18233 1847 18291 1853
rect 19334 1844 19340 1856
rect 19392 1844 19398 1896
rect 19705 1887 19763 1893
rect 19705 1853 19717 1887
rect 19751 1884 19763 1887
rect 19981 1887 20039 1893
rect 19751 1856 19932 1884
rect 19751 1853 19763 1856
rect 19705 1847 19763 1853
rect 19904 1748 19932 1856
rect 19981 1853 19993 1887
rect 20027 1853 20039 1887
rect 19981 1847 20039 1853
rect 19996 1816 20024 1847
rect 23198 1844 23204 1896
rect 23256 1844 23262 1896
rect 23569 1887 23627 1893
rect 23569 1853 23581 1887
rect 23615 1884 23627 1887
rect 24670 1884 24676 1896
rect 23615 1856 24676 1884
rect 23615 1853 23627 1856
rect 23569 1847 23627 1853
rect 24670 1844 24676 1856
rect 24728 1844 24734 1896
rect 25409 1887 25467 1893
rect 25409 1853 25421 1887
rect 25455 1884 25467 1887
rect 28442 1884 28448 1896
rect 25455 1856 28448 1884
rect 25455 1853 25467 1856
rect 25409 1847 25467 1853
rect 28442 1844 28448 1856
rect 28500 1844 28506 1896
rect 28721 1887 28779 1893
rect 28721 1853 28733 1887
rect 28767 1884 28779 1887
rect 28810 1884 28816 1896
rect 28767 1856 28816 1884
rect 28767 1853 28779 1856
rect 28721 1847 28779 1853
rect 28810 1844 28816 1856
rect 28868 1844 28874 1896
rect 28920 1884 28948 1915
rect 29086 1912 29092 1964
rect 29144 1912 29150 1964
rect 29546 1912 29552 1964
rect 29604 1952 29610 1964
rect 29748 1961 29776 1992
rect 66898 1980 66904 2032
rect 66956 2020 66962 2032
rect 66993 2023 67051 2029
rect 66993 2020 67005 2023
rect 66956 1992 67005 2020
rect 66956 1980 66962 1992
rect 66993 1989 67005 1992
rect 67039 1989 67051 2023
rect 67100 2020 67128 2060
rect 67266 2048 67272 2100
rect 67324 2048 67330 2100
rect 67910 2020 67916 2032
rect 67100 1992 67916 2020
rect 66993 1983 67051 1989
rect 67910 1980 67916 1992
rect 67968 1980 67974 2032
rect 69109 2023 69167 2029
rect 69109 1989 69121 2023
rect 69155 2020 69167 2023
rect 69198 2020 69204 2032
rect 69155 1992 69204 2020
rect 69155 1989 69167 1992
rect 69109 1983 69167 1989
rect 69198 1980 69204 1992
rect 69256 1980 69262 2032
rect 70118 1980 70124 2032
rect 70176 2020 70182 2032
rect 71961 2023 72019 2029
rect 71961 2020 71973 2023
rect 70176 1992 71973 2020
rect 70176 1980 70182 1992
rect 71961 1989 71973 1992
rect 72007 1989 72019 2023
rect 71961 1983 72019 1989
rect 29641 1955 29699 1961
rect 29641 1952 29653 1955
rect 29604 1924 29653 1952
rect 29604 1912 29610 1924
rect 29641 1921 29653 1924
rect 29687 1921 29699 1955
rect 29641 1915 29699 1921
rect 29733 1955 29791 1961
rect 29733 1921 29745 1955
rect 29779 1921 29791 1955
rect 29733 1915 29791 1921
rect 29914 1912 29920 1964
rect 29972 1952 29978 1964
rect 29972 1924 30420 1952
rect 29972 1912 29978 1924
rect 30282 1884 30288 1896
rect 28920 1856 30288 1884
rect 30282 1844 30288 1856
rect 30340 1844 30346 1896
rect 30392 1893 30420 1924
rect 31294 1912 31300 1964
rect 31352 1912 31358 1964
rect 33321 1955 33379 1961
rect 33321 1921 33333 1955
rect 33367 1952 33379 1955
rect 34054 1952 34060 1964
rect 33367 1924 34060 1952
rect 33367 1921 33379 1924
rect 33321 1915 33379 1921
rect 34054 1912 34060 1924
rect 34112 1912 34118 1964
rect 34790 1912 34796 1964
rect 34848 1912 34854 1964
rect 38105 1955 38163 1961
rect 38105 1921 38117 1955
rect 38151 1952 38163 1955
rect 38289 1955 38347 1961
rect 38289 1952 38301 1955
rect 38151 1924 38301 1952
rect 38151 1921 38163 1924
rect 38105 1915 38163 1921
rect 38289 1921 38301 1924
rect 38335 1921 38347 1955
rect 38289 1915 38347 1921
rect 39022 1912 39028 1964
rect 39080 1952 39086 1964
rect 40405 1955 40463 1961
rect 40405 1952 40417 1955
rect 39080 1924 40417 1952
rect 39080 1912 39086 1924
rect 40405 1921 40417 1924
rect 40451 1921 40463 1955
rect 40405 1915 40463 1921
rect 41693 1955 41751 1961
rect 41693 1921 41705 1955
rect 41739 1952 41751 1955
rect 41785 1955 41843 1961
rect 41785 1952 41797 1955
rect 41739 1924 41797 1952
rect 41739 1921 41751 1924
rect 41693 1915 41751 1921
rect 41785 1921 41797 1924
rect 41831 1921 41843 1955
rect 41785 1915 41843 1921
rect 42705 1955 42763 1961
rect 42705 1921 42717 1955
rect 42751 1952 42763 1955
rect 42886 1952 42892 1964
rect 42751 1924 42892 1952
rect 42751 1921 42763 1924
rect 42705 1915 42763 1921
rect 42886 1912 42892 1924
rect 42944 1912 42950 1964
rect 42978 1912 42984 1964
rect 43036 1912 43042 1964
rect 44729 1955 44787 1961
rect 44729 1921 44741 1955
rect 44775 1921 44787 1955
rect 44729 1915 44787 1921
rect 45373 1955 45431 1961
rect 45373 1921 45385 1955
rect 45419 1952 45431 1955
rect 45419 1924 45600 1952
rect 45419 1921 45431 1924
rect 45373 1915 45431 1921
rect 30377 1887 30435 1893
rect 30377 1853 30389 1887
rect 30423 1853 30435 1887
rect 30377 1847 30435 1853
rect 32398 1844 32404 1896
rect 32456 1884 32462 1896
rect 33137 1887 33195 1893
rect 33137 1884 33149 1887
rect 32456 1856 33149 1884
rect 32456 1844 32462 1856
rect 33137 1853 33149 1856
rect 33183 1853 33195 1887
rect 33137 1847 33195 1853
rect 33873 1887 33931 1893
rect 33873 1853 33885 1887
rect 33919 1884 33931 1887
rect 33965 1887 34023 1893
rect 33965 1884 33977 1887
rect 33919 1856 33977 1884
rect 33919 1853 33931 1856
rect 33873 1847 33931 1853
rect 33965 1853 33977 1856
rect 34011 1853 34023 1887
rect 33965 1847 34023 1853
rect 34606 1844 34612 1896
rect 34664 1884 34670 1896
rect 35161 1887 35219 1893
rect 35161 1884 35173 1887
rect 34664 1856 35173 1884
rect 34664 1844 34670 1856
rect 35161 1853 35173 1856
rect 35207 1853 35219 1887
rect 35161 1847 35219 1853
rect 36170 1844 36176 1896
rect 36228 1844 36234 1896
rect 37550 1844 37556 1896
rect 37608 1844 37614 1896
rect 39761 1887 39819 1893
rect 39761 1853 39773 1887
rect 39807 1884 39819 1887
rect 39853 1887 39911 1893
rect 39853 1884 39865 1887
rect 39807 1856 39865 1884
rect 39807 1853 39819 1856
rect 39761 1847 39819 1853
rect 39853 1853 39865 1856
rect 39899 1853 39911 1887
rect 39853 1847 39911 1853
rect 41138 1844 41144 1896
rect 41196 1844 41202 1896
rect 43441 1887 43499 1893
rect 43441 1853 43453 1887
rect 43487 1853 43499 1887
rect 44744 1884 44772 1915
rect 45465 1887 45523 1893
rect 45465 1884 45477 1887
rect 44744 1856 45477 1884
rect 43441 1847 43499 1853
rect 45465 1853 45477 1856
rect 45511 1853 45523 1887
rect 45465 1847 45523 1853
rect 35894 1816 35900 1828
rect 19996 1788 35900 1816
rect 35894 1776 35900 1788
rect 35952 1776 35958 1828
rect 35986 1776 35992 1828
rect 36044 1816 36050 1828
rect 41506 1816 41512 1828
rect 36044 1788 41512 1816
rect 36044 1776 36050 1788
rect 41506 1776 41512 1788
rect 41564 1776 41570 1828
rect 42978 1776 42984 1828
rect 43036 1816 43042 1828
rect 43456 1816 43484 1847
rect 43036 1788 43484 1816
rect 45572 1816 45600 1924
rect 45646 1912 45652 1964
rect 45704 1952 45710 1964
rect 46753 1955 46811 1961
rect 46753 1952 46765 1955
rect 45704 1924 46765 1952
rect 45704 1912 45710 1924
rect 46753 1921 46765 1924
rect 46799 1921 46811 1955
rect 46753 1915 46811 1921
rect 46842 1912 46848 1964
rect 46900 1952 46906 1964
rect 46937 1955 46995 1961
rect 46937 1952 46949 1955
rect 46900 1924 46949 1952
rect 46900 1912 46906 1924
rect 46937 1921 46949 1924
rect 46983 1921 46995 1955
rect 46937 1915 46995 1921
rect 47578 1912 47584 1964
rect 47636 1952 47642 1964
rect 47949 1955 48007 1961
rect 47949 1952 47961 1955
rect 47636 1924 47961 1952
rect 47636 1912 47642 1924
rect 47949 1921 47961 1924
rect 47995 1921 48007 1955
rect 47949 1915 48007 1921
rect 49510 1912 49516 1964
rect 49568 1912 49574 1964
rect 50065 1955 50123 1961
rect 50065 1921 50077 1955
rect 50111 1952 50123 1955
rect 50249 1955 50307 1961
rect 50249 1952 50261 1955
rect 50111 1924 50261 1952
rect 50111 1921 50123 1924
rect 50065 1915 50123 1921
rect 50249 1921 50261 1924
rect 50295 1921 50307 1955
rect 50249 1915 50307 1921
rect 51813 1955 51871 1961
rect 51813 1921 51825 1955
rect 51859 1952 51871 1955
rect 51997 1955 52055 1961
rect 51997 1952 52009 1955
rect 51859 1924 52009 1952
rect 51859 1921 51871 1924
rect 51813 1915 51871 1921
rect 51997 1921 52009 1924
rect 52043 1921 52055 1955
rect 51997 1915 52055 1921
rect 53098 1912 53104 1964
rect 53156 1912 53162 1964
rect 54481 1955 54539 1961
rect 54481 1921 54493 1955
rect 54527 1952 54539 1955
rect 54754 1952 54760 1964
rect 54527 1924 54760 1952
rect 54527 1921 54539 1924
rect 54481 1915 54539 1921
rect 54754 1912 54760 1924
rect 54812 1912 54818 1964
rect 56410 1912 56416 1964
rect 56468 1912 56474 1964
rect 57882 1912 57888 1964
rect 57940 1912 57946 1964
rect 58437 1955 58495 1961
rect 58437 1921 58449 1955
rect 58483 1952 58495 1955
rect 58621 1955 58679 1961
rect 58621 1952 58633 1955
rect 58483 1924 58633 1952
rect 58483 1921 58495 1924
rect 58437 1915 58495 1921
rect 58621 1921 58633 1924
rect 58667 1921 58679 1955
rect 58621 1915 58679 1921
rect 59817 1955 59875 1961
rect 59817 1921 59829 1955
rect 59863 1952 59875 1955
rect 60001 1955 60059 1961
rect 60001 1952 60013 1955
rect 59863 1924 60013 1952
rect 59863 1921 59875 1924
rect 59817 1915 59875 1921
rect 60001 1921 60013 1924
rect 60047 1921 60059 1955
rect 60001 1915 60059 1921
rect 61378 1912 61384 1964
rect 61436 1912 61442 1964
rect 62942 1912 62948 1964
rect 63000 1912 63006 1964
rect 64598 1912 64604 1964
rect 64656 1912 64662 1964
rect 66070 1912 66076 1964
rect 66128 1912 66134 1964
rect 66625 1955 66683 1961
rect 66625 1921 66637 1955
rect 66671 1952 66683 1955
rect 66717 1955 66775 1961
rect 66717 1952 66729 1955
rect 66671 1924 66729 1952
rect 66671 1921 66683 1924
rect 66625 1915 66683 1921
rect 66717 1921 66729 1924
rect 66763 1921 66775 1955
rect 66717 1915 66775 1921
rect 67174 1912 67180 1964
rect 67232 1952 67238 1964
rect 68649 1955 68707 1961
rect 68649 1952 68661 1955
rect 67232 1924 68661 1952
rect 67232 1912 67238 1924
rect 68649 1921 68661 1924
rect 68695 1921 68707 1955
rect 68649 1915 68707 1921
rect 69382 1912 69388 1964
rect 69440 1912 69446 1964
rect 69658 1912 69664 1964
rect 69716 1912 69722 1964
rect 71038 1912 71044 1964
rect 71096 1912 71102 1964
rect 71593 1955 71651 1961
rect 71593 1921 71605 1955
rect 71639 1952 71651 1955
rect 71685 1955 71743 1961
rect 71685 1952 71697 1955
rect 71639 1924 71697 1952
rect 71639 1921 71651 1924
rect 71593 1915 71651 1921
rect 71685 1921 71697 1924
rect 71731 1921 71743 1955
rect 71685 1915 71743 1921
rect 46014 1844 46020 1896
rect 46072 1844 46078 1896
rect 46198 1844 46204 1896
rect 46256 1844 46262 1896
rect 47854 1844 47860 1896
rect 47912 1884 47918 1896
rect 48409 1887 48467 1893
rect 48409 1884 48421 1887
rect 47912 1856 48421 1884
rect 47912 1844 47918 1856
rect 48409 1853 48421 1856
rect 48455 1853 48467 1887
rect 48409 1847 48467 1853
rect 51258 1844 51264 1896
rect 51316 1844 51322 1896
rect 52822 1844 52828 1896
rect 52880 1884 52886 1896
rect 53377 1887 53435 1893
rect 53377 1884 53389 1887
rect 52880 1856 53389 1884
rect 52880 1844 52886 1856
rect 53377 1853 53389 1856
rect 53423 1853 53435 1887
rect 53377 1847 53435 1853
rect 55582 1844 55588 1896
rect 55640 1844 55646 1896
rect 56134 1844 56140 1896
rect 56192 1884 56198 1896
rect 56689 1887 56747 1893
rect 56689 1884 56701 1887
rect 56192 1856 56701 1884
rect 56192 1844 56198 1856
rect 56689 1853 56701 1856
rect 56735 1853 56747 1887
rect 56689 1847 56747 1853
rect 59265 1887 59323 1893
rect 59265 1853 59277 1887
rect 59311 1884 59323 1887
rect 59354 1884 59360 1896
rect 59311 1856 59360 1884
rect 59311 1853 59323 1856
rect 59265 1847 59323 1853
rect 59354 1844 59360 1856
rect 59412 1844 59418 1896
rect 60550 1844 60556 1896
rect 60608 1844 60614 1896
rect 61102 1844 61108 1896
rect 61160 1884 61166 1896
rect 61657 1887 61715 1893
rect 61657 1884 61669 1887
rect 61160 1856 61669 1884
rect 61160 1844 61166 1856
rect 61657 1853 61669 1856
rect 61703 1853 61715 1887
rect 61657 1847 61715 1853
rect 63862 1844 63868 1896
rect 63920 1844 63926 1896
rect 64690 1844 64696 1896
rect 64748 1884 64754 1896
rect 64969 1887 65027 1893
rect 64969 1884 64981 1887
rect 64748 1856 64981 1884
rect 64748 1844 64754 1856
rect 64969 1853 64981 1856
rect 65015 1853 65027 1887
rect 64969 1847 65027 1853
rect 67913 1887 67971 1893
rect 67913 1853 67925 1887
rect 67959 1884 67971 1887
rect 68097 1887 68155 1893
rect 68097 1884 68109 1887
rect 67959 1856 68109 1884
rect 67959 1853 67971 1856
rect 67913 1847 67971 1853
rect 68097 1853 68109 1856
rect 68143 1853 68155 1887
rect 69937 1887 69995 1893
rect 69937 1884 69949 1887
rect 68097 1847 68155 1853
rect 69400 1856 69949 1884
rect 69400 1828 69428 1856
rect 69937 1853 69949 1856
rect 69983 1853 69995 1887
rect 69937 1847 69995 1853
rect 72234 1844 72240 1896
rect 72292 1884 72298 1896
rect 72329 1887 72387 1893
rect 72329 1884 72341 1887
rect 72292 1856 72341 1884
rect 72292 1844 72298 1856
rect 72329 1853 72341 1856
rect 72375 1853 72387 1887
rect 72329 1847 72387 1853
rect 72973 1887 73031 1893
rect 72973 1853 72985 1887
rect 73019 1884 73031 1887
rect 73801 1887 73859 1893
rect 73801 1884 73813 1887
rect 73019 1856 73813 1884
rect 73019 1853 73031 1856
rect 72973 1847 73031 1853
rect 73801 1853 73813 1856
rect 73847 1853 73859 1887
rect 73801 1847 73859 1853
rect 46934 1816 46940 1828
rect 45572 1788 46940 1816
rect 43036 1776 43042 1788
rect 46934 1776 46940 1788
rect 46992 1776 46998 1828
rect 52273 1819 52331 1825
rect 47044 1788 51074 1816
rect 23382 1748 23388 1760
rect 19904 1720 23388 1748
rect 23382 1708 23388 1720
rect 23440 1708 23446 1760
rect 28994 1708 29000 1760
rect 29052 1748 29058 1760
rect 34698 1748 34704 1760
rect 29052 1720 34704 1748
rect 29052 1708 29058 1720
rect 34698 1708 34704 1720
rect 34756 1708 34762 1760
rect 38562 1708 38568 1760
rect 38620 1708 38626 1760
rect 42521 1751 42579 1757
rect 42521 1717 42533 1751
rect 42567 1748 42579 1751
rect 47044 1748 47072 1788
rect 42567 1720 47072 1748
rect 47121 1751 47179 1757
rect 42567 1717 42579 1720
rect 42521 1711 42579 1717
rect 47121 1717 47133 1751
rect 47167 1748 47179 1751
rect 47210 1748 47216 1760
rect 47167 1720 47216 1748
rect 47167 1717 47179 1720
rect 47121 1711 47179 1717
rect 47210 1708 47216 1720
rect 47268 1708 47274 1760
rect 51046 1748 51074 1788
rect 52273 1785 52285 1819
rect 52319 1816 52331 1819
rect 55766 1816 55772 1828
rect 52319 1788 55772 1816
rect 52319 1785 52331 1788
rect 52273 1779 52331 1785
rect 55766 1776 55772 1788
rect 55824 1776 55830 1828
rect 60277 1819 60335 1825
rect 60277 1785 60289 1819
rect 60323 1816 60335 1819
rect 65426 1816 65432 1828
rect 60323 1788 65432 1816
rect 60323 1785 60335 1788
rect 60277 1779 60335 1785
rect 65426 1776 65432 1788
rect 65484 1776 65490 1828
rect 69382 1776 69388 1828
rect 69440 1776 69446 1828
rect 53374 1748 53380 1760
rect 51046 1720 53380 1748
rect 53374 1708 53380 1720
rect 53432 1708 53438 1760
rect 56137 1751 56195 1757
rect 56137 1717 56149 1751
rect 56183 1748 56195 1751
rect 57238 1748 57244 1760
rect 56183 1720 57244 1748
rect 56183 1717 56195 1720
rect 56137 1711 56195 1717
rect 57238 1708 57244 1720
rect 57296 1708 57302 1760
rect 61105 1751 61163 1757
rect 61105 1717 61117 1751
rect 61151 1748 61163 1751
rect 62390 1748 62396 1760
rect 61151 1720 62396 1748
rect 61151 1717 61163 1720
rect 61105 1711 61163 1717
rect 62390 1708 62396 1720
rect 62448 1708 62454 1760
rect 64417 1751 64475 1757
rect 64417 1717 64429 1751
rect 64463 1748 64475 1751
rect 65150 1748 65156 1760
rect 64463 1720 65156 1748
rect 64463 1717 64475 1720
rect 64417 1711 64475 1717
rect 65150 1708 65156 1720
rect 65208 1708 65214 1760
rect 73154 1708 73160 1760
rect 73212 1748 73218 1760
rect 73249 1751 73307 1757
rect 73249 1748 73261 1751
rect 73212 1720 73261 1748
rect 73212 1708 73218 1720
rect 73249 1717 73261 1720
rect 73295 1717 73307 1751
rect 73249 1711 73307 1717
rect 1012 1658 74980 1680
rect 1012 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 74980 1658
rect 1012 1584 74980 1606
rect 22649 1547 22707 1553
rect 22649 1513 22661 1547
rect 22695 1544 22707 1547
rect 22922 1544 22928 1556
rect 22695 1516 22928 1544
rect 22695 1513 22707 1516
rect 22649 1507 22707 1513
rect 22922 1504 22928 1516
rect 22980 1504 22986 1556
rect 25225 1547 25283 1553
rect 25225 1513 25237 1547
rect 25271 1544 25283 1547
rect 26050 1544 26056 1556
rect 25271 1516 26056 1544
rect 25271 1513 25283 1516
rect 25225 1507 25283 1513
rect 26050 1504 26056 1516
rect 26108 1504 26114 1556
rect 27801 1547 27859 1553
rect 27801 1513 27813 1547
rect 27847 1544 27859 1547
rect 28626 1544 28632 1556
rect 27847 1516 28632 1544
rect 27847 1513 27859 1516
rect 27801 1507 27859 1513
rect 28626 1504 28632 1516
rect 28684 1504 28690 1556
rect 30377 1547 30435 1553
rect 30377 1513 30389 1547
rect 30423 1544 30435 1547
rect 31018 1544 31024 1556
rect 30423 1516 31024 1544
rect 30423 1513 30435 1516
rect 30377 1507 30435 1513
rect 31018 1504 31024 1516
rect 31076 1504 31082 1556
rect 37550 1504 37556 1556
rect 37608 1544 37614 1556
rect 37921 1547 37979 1553
rect 37921 1544 37933 1547
rect 37608 1516 37933 1544
rect 37608 1504 37614 1516
rect 37921 1513 37933 1516
rect 37967 1513 37979 1547
rect 37921 1507 37979 1513
rect 41138 1504 41144 1556
rect 41196 1544 41202 1556
rect 41233 1547 41291 1553
rect 41233 1544 41245 1547
rect 41196 1516 41245 1544
rect 41196 1504 41202 1516
rect 41233 1513 41245 1516
rect 41279 1513 41291 1547
rect 45462 1544 45468 1556
rect 41233 1507 41291 1513
rect 41386 1516 45468 1544
rect 31110 1476 31116 1488
rect 22066 1448 31116 1476
rect 20993 1411 21051 1417
rect 20993 1377 21005 1411
rect 21039 1408 21051 1411
rect 22066 1408 22094 1448
rect 31110 1436 31116 1448
rect 31168 1436 31174 1488
rect 35158 1436 35164 1488
rect 35216 1476 35222 1488
rect 36538 1476 36544 1488
rect 35216 1448 36544 1476
rect 35216 1436 35222 1448
rect 36538 1436 36544 1448
rect 36596 1436 36602 1488
rect 38562 1436 38568 1488
rect 38620 1476 38626 1488
rect 41386 1476 41414 1516
rect 45462 1504 45468 1516
rect 45520 1504 45526 1556
rect 45554 1504 45560 1556
rect 45612 1544 45618 1556
rect 46385 1547 46443 1553
rect 46385 1544 46397 1547
rect 45612 1516 46397 1544
rect 45612 1504 45618 1516
rect 46385 1513 46397 1516
rect 46431 1513 46443 1547
rect 46385 1507 46443 1513
rect 46934 1504 46940 1556
rect 46992 1544 46998 1556
rect 47121 1547 47179 1553
rect 47121 1544 47133 1547
rect 46992 1516 47133 1544
rect 46992 1504 46998 1516
rect 47121 1513 47133 1516
rect 47167 1513 47179 1547
rect 47121 1507 47179 1513
rect 51258 1504 51264 1556
rect 51316 1544 51322 1556
rect 51537 1547 51595 1553
rect 51537 1544 51549 1547
rect 51316 1516 51549 1544
rect 51316 1504 51322 1516
rect 51537 1513 51549 1516
rect 51583 1513 51595 1547
rect 51537 1507 51595 1513
rect 61010 1504 61016 1556
rect 61068 1544 61074 1556
rect 61841 1547 61899 1553
rect 61841 1544 61853 1547
rect 61068 1516 61853 1544
rect 61068 1504 61074 1516
rect 61841 1513 61853 1516
rect 61887 1513 61899 1547
rect 61841 1507 61899 1513
rect 63862 1504 63868 1556
rect 63920 1544 63926 1556
rect 64417 1547 64475 1553
rect 64417 1544 64429 1547
rect 63920 1516 64429 1544
rect 63920 1504 63926 1516
rect 64417 1513 64429 1516
rect 64463 1513 64475 1547
rect 64417 1507 64475 1513
rect 69934 1504 69940 1556
rect 69992 1544 69998 1556
rect 70213 1547 70271 1553
rect 70213 1544 70225 1547
rect 69992 1516 70225 1544
rect 69992 1504 69998 1516
rect 70213 1513 70225 1516
rect 70259 1513 70271 1547
rect 70213 1507 70271 1513
rect 38620 1448 41414 1476
rect 38620 1436 38626 1448
rect 41690 1436 41696 1488
rect 41748 1476 41754 1488
rect 47026 1476 47032 1488
rect 41748 1448 47032 1476
rect 41748 1436 41754 1448
rect 47026 1436 47032 1448
rect 47084 1436 47090 1488
rect 21039 1380 22094 1408
rect 21039 1377 21051 1380
rect 20993 1371 21051 1377
rect 27982 1368 27988 1420
rect 28040 1408 28046 1420
rect 28353 1411 28411 1417
rect 28353 1408 28365 1411
rect 28040 1380 28365 1408
rect 28040 1368 28046 1380
rect 28353 1377 28365 1380
rect 28399 1377 28411 1411
rect 28353 1371 28411 1377
rect 28442 1368 28448 1420
rect 28500 1408 28506 1420
rect 35066 1408 35072 1420
rect 28500 1380 35072 1408
rect 28500 1368 28506 1380
rect 35066 1368 35072 1380
rect 35124 1368 35130 1420
rect 37918 1368 37924 1420
rect 37976 1408 37982 1420
rect 38473 1411 38531 1417
rect 38473 1408 38485 1411
rect 37976 1380 38485 1408
rect 37976 1368 37982 1380
rect 38473 1377 38485 1380
rect 38519 1377 38531 1411
rect 38473 1371 38531 1377
rect 41230 1368 41236 1420
rect 41288 1408 41294 1420
rect 42797 1411 42855 1417
rect 42797 1408 42809 1411
rect 41288 1380 42809 1408
rect 41288 1368 41294 1380
rect 42797 1377 42809 1380
rect 42843 1377 42855 1411
rect 44634 1408 44640 1420
rect 42797 1371 42855 1377
rect 44468 1380 44640 1408
rect 5074 1300 5080 1352
rect 5132 1300 5138 1352
rect 15286 1300 15292 1352
rect 15344 1340 15350 1352
rect 15381 1343 15439 1349
rect 15381 1340 15393 1343
rect 15344 1312 15393 1340
rect 15344 1300 15350 1312
rect 15381 1309 15393 1312
rect 15427 1309 15439 1343
rect 15381 1303 15439 1309
rect 15841 1343 15899 1349
rect 15841 1309 15853 1343
rect 15887 1340 15899 1343
rect 17494 1340 17500 1352
rect 15887 1312 17500 1340
rect 15887 1309 15899 1312
rect 15841 1303 15899 1309
rect 17494 1300 17500 1312
rect 17552 1300 17558 1352
rect 17770 1300 17776 1352
rect 17828 1300 17834 1352
rect 18049 1343 18107 1349
rect 18049 1309 18061 1343
rect 18095 1309 18107 1343
rect 18049 1303 18107 1309
rect 18325 1343 18383 1349
rect 18325 1309 18337 1343
rect 18371 1340 18383 1343
rect 19058 1340 19064 1352
rect 18371 1312 19064 1340
rect 18371 1309 18383 1312
rect 18325 1303 18383 1309
rect 3142 1232 3148 1284
rect 3200 1272 3206 1284
rect 3881 1275 3939 1281
rect 3881 1272 3893 1275
rect 3200 1244 3893 1272
rect 3200 1232 3206 1244
rect 3881 1241 3893 1244
rect 3927 1241 3939 1275
rect 3881 1235 3939 1241
rect 15930 1232 15936 1284
rect 15988 1272 15994 1284
rect 16761 1275 16819 1281
rect 16761 1272 16773 1275
rect 15988 1244 16773 1272
rect 15988 1232 15994 1244
rect 16761 1241 16773 1244
rect 16807 1241 16819 1275
rect 16761 1235 16819 1241
rect 15562 1164 15568 1216
rect 15620 1164 15626 1216
rect 16393 1207 16451 1213
rect 16393 1173 16405 1207
rect 16439 1204 16451 1207
rect 18064 1204 18092 1303
rect 19058 1300 19064 1312
rect 19116 1300 19122 1352
rect 19705 1343 19763 1349
rect 19705 1309 19717 1343
rect 19751 1309 19763 1343
rect 19705 1303 19763 1309
rect 19426 1232 19432 1284
rect 19484 1232 19490 1284
rect 19720 1272 19748 1303
rect 19794 1300 19800 1352
rect 19852 1300 19858 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22554 1340 22560 1352
rect 22051 1312 22560 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22554 1300 22560 1312
rect 22612 1300 22618 1352
rect 24121 1343 24179 1349
rect 24121 1309 24133 1343
rect 24167 1309 24179 1343
rect 24121 1303 24179 1309
rect 24673 1343 24731 1349
rect 24673 1309 24685 1343
rect 24719 1340 24731 1343
rect 26326 1340 26332 1352
rect 24719 1312 26332 1340
rect 24719 1309 24731 1312
rect 24673 1303 24731 1309
rect 22278 1272 22284 1284
rect 19720 1244 22284 1272
rect 22278 1232 22284 1244
rect 22336 1232 22342 1284
rect 23201 1275 23259 1281
rect 23201 1241 23213 1275
rect 23247 1272 23259 1275
rect 23566 1272 23572 1284
rect 23247 1244 23572 1272
rect 23247 1241 23259 1244
rect 23201 1235 23259 1241
rect 23566 1232 23572 1244
rect 23624 1232 23630 1284
rect 16439 1176 18092 1204
rect 24136 1204 24164 1303
rect 26326 1300 26332 1312
rect 26384 1300 26390 1352
rect 26697 1343 26755 1349
rect 26697 1309 26709 1343
rect 26743 1309 26755 1343
rect 26697 1303 26755 1309
rect 27249 1343 27307 1349
rect 27249 1309 27261 1343
rect 27295 1309 27307 1343
rect 27249 1303 27307 1309
rect 25774 1232 25780 1284
rect 25832 1232 25838 1284
rect 26510 1204 26516 1216
rect 24136 1176 26516 1204
rect 16439 1173 16451 1176
rect 16393 1167 16451 1173
rect 26510 1164 26516 1176
rect 26568 1164 26574 1216
rect 26712 1204 26740 1303
rect 27264 1272 27292 1303
rect 28074 1300 28080 1352
rect 28132 1300 28138 1352
rect 29454 1300 29460 1352
rect 29512 1300 29518 1352
rect 29825 1343 29883 1349
rect 29825 1309 29837 1343
rect 29871 1340 29883 1343
rect 30374 1340 30380 1352
rect 29871 1312 30380 1340
rect 29871 1309 29883 1312
rect 29825 1303 29883 1309
rect 30374 1300 30380 1312
rect 30432 1300 30438 1352
rect 30469 1343 30527 1349
rect 30469 1309 30481 1343
rect 30515 1309 30527 1343
rect 30469 1303 30527 1309
rect 32401 1343 32459 1349
rect 32401 1309 32413 1343
rect 32447 1340 32459 1343
rect 32858 1340 32864 1352
rect 32447 1312 32864 1340
rect 32447 1309 32459 1312
rect 32401 1303 32459 1309
rect 28534 1272 28540 1284
rect 27264 1244 28540 1272
rect 28534 1232 28540 1244
rect 28592 1232 28598 1284
rect 30484 1272 30512 1303
rect 32858 1300 32864 1312
rect 32916 1300 32922 1352
rect 33226 1300 33232 1352
rect 33284 1300 33290 1352
rect 34977 1343 35035 1349
rect 34977 1309 34989 1343
rect 35023 1309 35035 1343
rect 34977 1303 35035 1309
rect 29656 1244 30512 1272
rect 27890 1204 27896 1216
rect 26712 1176 27896 1204
rect 27890 1164 27896 1176
rect 27948 1164 27954 1216
rect 29656 1213 29684 1244
rect 31294 1232 31300 1284
rect 31352 1272 31358 1284
rect 31389 1275 31447 1281
rect 31389 1272 31401 1275
rect 31352 1244 31401 1272
rect 31352 1232 31358 1244
rect 31389 1241 31401 1244
rect 31435 1241 31447 1275
rect 31389 1235 31447 1241
rect 33042 1232 33048 1284
rect 33100 1272 33106 1284
rect 33965 1275 34023 1281
rect 33965 1272 33977 1275
rect 33100 1244 33977 1272
rect 33100 1232 33106 1244
rect 33965 1241 33977 1244
rect 34011 1241 34023 1275
rect 33965 1235 34023 1241
rect 29641 1207 29699 1213
rect 29641 1173 29653 1207
rect 29687 1173 29699 1207
rect 29641 1167 29699 1173
rect 32953 1207 33011 1213
rect 32953 1173 32965 1207
rect 32999 1204 33011 1207
rect 33594 1204 33600 1216
rect 32999 1176 33600 1204
rect 32999 1173 33011 1176
rect 32953 1167 33011 1173
rect 33594 1164 33600 1176
rect 33652 1164 33658 1216
rect 34992 1204 35020 1303
rect 35618 1300 35624 1352
rect 35676 1300 35682 1352
rect 37366 1300 37372 1352
rect 37424 1300 37430 1352
rect 38010 1300 38016 1352
rect 38068 1300 38074 1352
rect 39758 1300 39764 1352
rect 39816 1300 39822 1352
rect 40770 1300 40776 1352
rect 40828 1340 40834 1352
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 40828 1312 41797 1340
rect 40828 1300 40834 1312
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41785 1303 41843 1309
rect 42426 1300 42432 1352
rect 42484 1300 42490 1352
rect 42886 1300 42892 1352
rect 42944 1340 42950 1352
rect 44468 1349 44496 1380
rect 44634 1368 44640 1380
rect 44692 1368 44698 1420
rect 44818 1368 44824 1420
rect 44876 1408 44882 1420
rect 45373 1411 45431 1417
rect 45373 1408 45385 1411
rect 44876 1380 45385 1408
rect 44876 1368 44882 1380
rect 45373 1377 45385 1380
rect 45419 1377 45431 1411
rect 45373 1371 45431 1377
rect 46198 1368 46204 1420
rect 46256 1408 46262 1420
rect 47949 1411 48007 1417
rect 47949 1408 47961 1411
rect 46256 1380 47961 1408
rect 46256 1368 46262 1380
rect 47949 1377 47961 1380
rect 47995 1377 48007 1411
rect 47949 1371 48007 1377
rect 49602 1368 49608 1420
rect 49660 1408 49666 1420
rect 50525 1411 50583 1417
rect 50525 1408 50537 1411
rect 49660 1380 50537 1408
rect 49660 1368 49666 1380
rect 50525 1377 50537 1380
rect 50571 1377 50583 1411
rect 50525 1371 50583 1377
rect 59446 1368 59452 1420
rect 59504 1408 59510 1420
rect 60829 1411 60887 1417
rect 60829 1408 60841 1411
rect 59504 1380 60841 1408
rect 59504 1368 59510 1380
rect 60829 1377 60841 1380
rect 60875 1377 60887 1411
rect 60829 1371 60887 1377
rect 62758 1368 62764 1420
rect 62816 1408 62822 1420
rect 63405 1411 63463 1417
rect 63405 1408 63417 1411
rect 62816 1380 63417 1408
rect 62816 1368 62822 1380
rect 63405 1377 63417 1380
rect 63451 1377 63463 1411
rect 63405 1371 63463 1377
rect 67726 1368 67732 1420
rect 67784 1408 67790 1420
rect 68557 1411 68615 1417
rect 68557 1408 68569 1411
rect 67784 1380 68569 1408
rect 67784 1368 67790 1380
rect 68557 1377 68569 1380
rect 68603 1377 68615 1411
rect 68557 1371 68615 1377
rect 71038 1368 71044 1420
rect 71096 1408 71102 1420
rect 71593 1411 71651 1417
rect 71593 1408 71605 1411
rect 71096 1380 71605 1408
rect 71096 1368 71102 1380
rect 71593 1377 71605 1380
rect 71639 1377 71651 1411
rect 71593 1371 71651 1377
rect 43809 1343 43867 1349
rect 43809 1340 43821 1343
rect 42944 1312 43821 1340
rect 42944 1300 42950 1312
rect 43809 1309 43821 1312
rect 43855 1309 43867 1343
rect 43809 1303 43867 1309
rect 44453 1343 44511 1349
rect 44453 1309 44465 1343
rect 44499 1309 44511 1343
rect 44453 1303 44511 1309
rect 44545 1343 44603 1349
rect 44545 1309 44557 1343
rect 44591 1340 44603 1343
rect 44726 1340 44732 1352
rect 44591 1312 44732 1340
rect 44591 1309 44603 1312
rect 44545 1303 44603 1309
rect 44726 1300 44732 1312
rect 44784 1300 44790 1352
rect 44910 1300 44916 1352
rect 44968 1300 44974 1352
rect 46937 1343 46995 1349
rect 46937 1340 46949 1343
rect 45020 1312 46949 1340
rect 35529 1275 35587 1281
rect 35529 1241 35541 1275
rect 35575 1272 35587 1275
rect 36170 1272 36176 1284
rect 35575 1244 36176 1272
rect 35575 1241 35587 1244
rect 35529 1235 35587 1241
rect 36170 1232 36176 1244
rect 36228 1232 36234 1284
rect 36262 1232 36268 1284
rect 36320 1272 36326 1284
rect 36541 1275 36599 1281
rect 36541 1272 36553 1275
rect 36320 1244 36553 1272
rect 36320 1232 36326 1244
rect 36541 1241 36553 1244
rect 36587 1241 36599 1275
rect 36541 1235 36599 1241
rect 39574 1232 39580 1284
rect 39632 1272 39638 1284
rect 40681 1275 40739 1281
rect 40681 1272 40693 1275
rect 39632 1244 40693 1272
rect 39632 1232 39638 1244
rect 40681 1241 40693 1244
rect 40727 1241 40739 1275
rect 40681 1235 40739 1241
rect 43990 1232 43996 1284
rect 44048 1272 44054 1284
rect 45020 1272 45048 1312
rect 46937 1309 46949 1312
rect 46983 1309 46995 1343
rect 46937 1303 46995 1309
rect 47305 1343 47363 1349
rect 47305 1309 47317 1343
rect 47351 1309 47363 1343
rect 47305 1303 47363 1309
rect 44048 1244 45048 1272
rect 44048 1232 44054 1244
rect 45094 1232 45100 1284
rect 45152 1272 45158 1284
rect 47320 1272 47348 1303
rect 47486 1300 47492 1352
rect 47544 1300 47550 1352
rect 48866 1300 48872 1352
rect 48924 1340 48930 1352
rect 48961 1343 49019 1349
rect 48961 1340 48973 1343
rect 48924 1312 48973 1340
rect 48924 1300 48930 1312
rect 48961 1309 48973 1312
rect 49007 1309 49019 1343
rect 48961 1303 49019 1309
rect 49418 1300 49424 1352
rect 49476 1340 49482 1352
rect 49513 1343 49571 1349
rect 49513 1340 49525 1343
rect 49476 1312 49525 1340
rect 49476 1300 49482 1312
rect 49513 1309 49525 1312
rect 49559 1309 49571 1343
rect 49513 1303 49571 1309
rect 50062 1300 50068 1352
rect 50120 1300 50126 1352
rect 50614 1300 50620 1352
rect 50672 1340 50678 1352
rect 52089 1343 52147 1349
rect 52089 1340 52101 1343
rect 50672 1312 52101 1340
rect 50672 1300 50678 1312
rect 52089 1309 52101 1312
rect 52135 1309 52147 1343
rect 52089 1303 52147 1309
rect 52638 1300 52644 1352
rect 52696 1300 52702 1352
rect 53834 1300 53840 1352
rect 53892 1340 53898 1352
rect 54113 1343 54171 1349
rect 54113 1340 54125 1343
rect 53892 1312 54125 1340
rect 53892 1300 53898 1312
rect 54113 1309 54125 1312
rect 54159 1309 54171 1343
rect 54665 1343 54723 1349
rect 54665 1340 54677 1343
rect 54113 1303 54171 1309
rect 54220 1312 54677 1340
rect 45152 1244 47348 1272
rect 45152 1232 45158 1244
rect 51166 1232 51172 1284
rect 51224 1272 51230 1284
rect 53561 1275 53619 1281
rect 53561 1272 53573 1275
rect 51224 1244 53573 1272
rect 51224 1232 51230 1244
rect 53561 1241 53573 1244
rect 53607 1241 53619 1275
rect 53561 1235 53619 1241
rect 35710 1204 35716 1216
rect 34992 1176 35716 1204
rect 35710 1164 35716 1176
rect 35768 1164 35774 1216
rect 44729 1207 44787 1213
rect 44729 1173 44741 1207
rect 44775 1204 44787 1207
rect 46014 1204 46020 1216
rect 44775 1176 46020 1204
rect 44775 1173 44787 1176
rect 44729 1167 44787 1173
rect 46014 1164 46020 1176
rect 46072 1164 46078 1216
rect 52270 1164 52276 1216
rect 52328 1204 52334 1216
rect 54220 1204 54248 1312
rect 54665 1309 54677 1312
rect 54711 1309 54723 1343
rect 54665 1303 54723 1309
rect 55214 1300 55220 1352
rect 55272 1300 55278 1352
rect 56686 1300 56692 1352
rect 56744 1300 56750 1352
rect 57238 1300 57244 1352
rect 57296 1300 57302 1352
rect 57974 1300 57980 1352
rect 58032 1300 58038 1352
rect 59354 1300 59360 1352
rect 59412 1300 59418 1352
rect 59909 1343 59967 1349
rect 59909 1309 59921 1343
rect 59955 1309 59967 1343
rect 59909 1303 59967 1309
rect 54570 1232 54576 1284
rect 54628 1272 54634 1284
rect 56137 1275 56195 1281
rect 56137 1272 56149 1275
rect 54628 1244 56149 1272
rect 54628 1232 54634 1244
rect 56137 1241 56149 1244
rect 56183 1241 56195 1275
rect 56137 1235 56195 1241
rect 57790 1232 57796 1284
rect 57848 1272 57854 1284
rect 58805 1275 58863 1281
rect 58805 1272 58817 1275
rect 57848 1244 58817 1272
rect 57848 1232 57854 1244
rect 58805 1241 58817 1244
rect 58851 1241 58863 1275
rect 58805 1235 58863 1241
rect 58894 1232 58900 1284
rect 58952 1272 58958 1284
rect 59924 1272 59952 1303
rect 60366 1300 60372 1352
rect 60424 1300 60430 1352
rect 62390 1300 62396 1352
rect 62448 1300 62454 1352
rect 63034 1300 63040 1352
rect 63092 1300 63098 1352
rect 63862 1300 63868 1352
rect 63920 1340 63926 1352
rect 64969 1343 65027 1349
rect 64969 1340 64981 1343
rect 63920 1312 64981 1340
rect 63920 1300 63926 1312
rect 64969 1309 64981 1312
rect 65015 1309 65027 1343
rect 64969 1303 65027 1309
rect 65150 1300 65156 1352
rect 65208 1340 65214 1352
rect 65521 1343 65579 1349
rect 65521 1340 65533 1343
rect 65208 1312 65533 1340
rect 65208 1300 65214 1312
rect 65521 1309 65533 1312
rect 65567 1309 65579 1343
rect 65521 1303 65579 1309
rect 66254 1300 66260 1352
rect 66312 1300 66318 1352
rect 68278 1300 68284 1352
rect 68336 1300 68342 1352
rect 68830 1300 68836 1352
rect 68888 1340 68894 1352
rect 69569 1343 69627 1349
rect 69569 1340 69581 1343
rect 68888 1312 69581 1340
rect 68888 1300 68894 1312
rect 69569 1309 69581 1312
rect 69615 1309 69627 1343
rect 69569 1303 69627 1309
rect 71222 1300 71228 1352
rect 71280 1300 71286 1352
rect 73065 1343 73123 1349
rect 73065 1309 73077 1343
rect 73111 1340 73123 1343
rect 73154 1340 73160 1352
rect 73111 1312 73160 1340
rect 73111 1309 73123 1312
rect 73065 1303 73123 1309
rect 73154 1300 73160 1312
rect 73212 1300 73218 1352
rect 73246 1300 73252 1352
rect 73304 1300 73310 1352
rect 58952 1244 59952 1272
rect 65797 1275 65855 1281
rect 58952 1232 58958 1244
rect 65797 1241 65809 1275
rect 65843 1241 65855 1275
rect 65797 1235 65855 1241
rect 52328 1176 54248 1204
rect 65812 1204 65840 1235
rect 66070 1232 66076 1284
rect 66128 1272 66134 1284
rect 67085 1275 67143 1281
rect 67085 1272 67097 1275
rect 66128 1244 67097 1272
rect 66128 1232 66134 1244
rect 67085 1241 67097 1244
rect 67131 1241 67143 1275
rect 67085 1235 67143 1241
rect 70026 1232 70032 1284
rect 70084 1272 70090 1284
rect 72789 1275 72847 1281
rect 72789 1272 72801 1275
rect 70084 1244 72801 1272
rect 70084 1232 70090 1244
rect 72789 1241 72801 1244
rect 72835 1241 72847 1275
rect 72789 1235 72847 1241
rect 74169 1275 74227 1281
rect 74169 1241 74181 1275
rect 74215 1241 74227 1275
rect 74169 1235 74227 1241
rect 67358 1204 67364 1216
rect 65812 1176 67364 1204
rect 52328 1164 52334 1176
rect 67358 1164 67364 1176
rect 67416 1164 67422 1216
rect 72694 1164 72700 1216
rect 72752 1204 72758 1216
rect 74184 1204 74212 1235
rect 72752 1176 74212 1204
rect 72752 1164 72758 1176
rect 1012 1114 74980 1136
rect 1012 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74980 1114
rect 1012 1040 74980 1062
rect 5074 960 5080 1012
rect 5132 1000 5138 1012
rect 23934 1000 23940 1012
rect 5132 972 23940 1000
rect 5132 960 5138 972
rect 23934 960 23940 972
rect 23992 960 23998 1012
rect 31386 960 31392 1012
rect 31444 1000 31450 1012
rect 35618 1000 35624 1012
rect 31444 972 35624 1000
rect 31444 960 31450 972
rect 35618 960 35624 972
rect 35676 960 35682 1012
rect 15562 892 15568 944
rect 15620 932 15626 944
rect 20714 932 20720 944
rect 15620 904 20720 932
rect 15620 892 15626 904
rect 20714 892 20720 904
rect 20772 892 20778 944
rect 32858 892 32864 944
rect 32916 932 32922 944
rect 33502 932 33508 944
rect 32916 904 33508 932
rect 32916 892 32922 904
rect 33502 892 33508 904
rect 33560 892 33566 944
rect 19426 824 19432 876
rect 19484 864 19490 876
rect 43806 864 43812 876
rect 19484 836 43812 864
rect 19484 824 19490 836
rect 43806 824 43812 836
rect 43864 824 43870 876
<< via1 >>
rect 74210 85926 74262 85978
rect 74274 85926 74326 85978
rect 74338 85926 74390 85978
rect 74402 85926 74454 85978
rect 74466 85926 74518 85978
rect 71858 85382 71910 85434
rect 71922 85382 71974 85434
rect 71986 85382 72038 85434
rect 72050 85382 72102 85434
rect 72114 85382 72166 85434
rect 74210 84838 74262 84890
rect 74274 84838 74326 84890
rect 74338 84838 74390 84890
rect 74402 84838 74454 84890
rect 74466 84838 74518 84890
rect 71858 84294 71910 84346
rect 71922 84294 71974 84346
rect 71986 84294 72038 84346
rect 72050 84294 72102 84346
rect 72114 84294 72166 84346
rect 64880 84192 64932 84244
rect 74210 83750 74262 83802
rect 74274 83750 74326 83802
rect 74338 83750 74390 83802
rect 74402 83750 74454 83802
rect 74466 83750 74518 83802
rect 71858 83206 71910 83258
rect 71922 83206 71974 83258
rect 71986 83206 72038 83258
rect 72050 83206 72102 83258
rect 72114 83206 72166 83258
rect 66996 83104 67048 83156
rect 69664 82968 69716 83020
rect 74210 82662 74262 82714
rect 74274 82662 74326 82714
rect 74338 82662 74390 82714
rect 74402 82662 74454 82714
rect 74466 82662 74518 82714
rect 71858 82118 71910 82170
rect 71922 82118 71974 82170
rect 71986 82118 72038 82170
rect 72050 82118 72102 82170
rect 72114 82118 72166 82170
rect 64880 81744 64932 81796
rect 74210 81574 74262 81626
rect 74274 81574 74326 81626
rect 74338 81574 74390 81626
rect 74402 81574 74454 81626
rect 74466 81574 74518 81626
rect 71858 81030 71910 81082
rect 71922 81030 71974 81082
rect 71986 81030 72038 81082
rect 72050 81030 72102 81082
rect 72114 81030 72166 81082
rect 67088 80928 67140 80980
rect 69756 80792 69808 80844
rect 74210 80486 74262 80538
rect 74274 80486 74326 80538
rect 74338 80486 74390 80538
rect 74402 80486 74454 80538
rect 74466 80486 74518 80538
rect 71858 79942 71910 79994
rect 71922 79942 71974 79994
rect 71986 79942 72038 79994
rect 72050 79942 72102 79994
rect 72114 79942 72166 79994
rect 64880 79840 64932 79892
rect 74210 79398 74262 79450
rect 74274 79398 74326 79450
rect 74338 79398 74390 79450
rect 74402 79398 74454 79450
rect 74466 79398 74518 79450
rect 71858 78854 71910 78906
rect 71922 78854 71974 78906
rect 71986 78854 72038 78906
rect 72050 78854 72102 78906
rect 72114 78854 72166 78906
rect 66444 78684 66496 78736
rect 69940 78616 69992 78668
rect 74210 78310 74262 78362
rect 74274 78310 74326 78362
rect 74338 78310 74390 78362
rect 74402 78310 74454 78362
rect 74466 78310 74518 78362
rect 71858 77766 71910 77818
rect 71922 77766 71974 77818
rect 71986 77766 72038 77818
rect 72050 77766 72102 77818
rect 72114 77766 72166 77818
rect 64880 77664 64932 77716
rect 74210 77222 74262 77274
rect 74274 77222 74326 77274
rect 74338 77222 74390 77274
rect 74402 77222 74454 77274
rect 74466 77222 74518 77274
rect 71858 76678 71910 76730
rect 71922 76678 71974 76730
rect 71986 76678 72038 76730
rect 72050 76678 72102 76730
rect 72114 76678 72166 76730
rect 66260 76508 66312 76560
rect 68468 76440 68520 76492
rect 74210 76134 74262 76186
rect 74274 76134 74326 76186
rect 74338 76134 74390 76186
rect 74402 76134 74454 76186
rect 74466 76134 74518 76186
rect 71858 75590 71910 75642
rect 71922 75590 71974 75642
rect 71986 75590 72038 75642
rect 72050 75590 72102 75642
rect 72114 75590 72166 75642
rect 64880 75148 64932 75200
rect 74210 75046 74262 75098
rect 74274 75046 74326 75098
rect 74338 75046 74390 75098
rect 74402 75046 74454 75098
rect 74466 75046 74518 75098
rect 67824 74604 67876 74656
rect 71858 74502 71910 74554
rect 71922 74502 71974 74554
rect 71986 74502 72038 74554
rect 72050 74502 72102 74554
rect 72114 74502 72166 74554
rect 66168 74060 66220 74112
rect 74210 73958 74262 74010
rect 74274 73958 74326 74010
rect 74338 73958 74390 74010
rect 74402 73958 74454 74010
rect 74466 73958 74518 74010
rect 71858 73414 71910 73466
rect 71922 73414 71974 73466
rect 71986 73414 72038 73466
rect 72050 73414 72102 73466
rect 72114 73414 72166 73466
rect 64880 73176 64932 73228
rect 74210 72870 74262 72922
rect 74274 72870 74326 72922
rect 74338 72870 74390 72922
rect 74402 72870 74454 72922
rect 74466 72870 74518 72922
rect 71858 72326 71910 72378
rect 71922 72326 71974 72378
rect 71986 72326 72038 72378
rect 72050 72326 72102 72378
rect 72114 72326 72166 72378
rect 66628 72156 66680 72208
rect 65064 71748 65116 71800
rect 74210 71782 74262 71834
rect 74274 71782 74326 71834
rect 74338 71782 74390 71834
rect 74402 71782 74454 71834
rect 74466 71782 74518 71834
rect 71858 71238 71910 71290
rect 71922 71238 71974 71290
rect 71986 71238 72038 71290
rect 72050 71238 72102 71290
rect 72114 71238 72166 71290
rect 64880 71068 64932 71120
rect 74210 70694 74262 70746
rect 74274 70694 74326 70746
rect 74338 70694 74390 70746
rect 74402 70694 74454 70746
rect 74466 70694 74518 70746
rect 71858 70150 71910 70202
rect 71922 70150 71974 70202
rect 71986 70150 72038 70202
rect 72050 70150 72102 70202
rect 72114 70150 72166 70202
rect 65524 69980 65576 70032
rect 63684 69572 63736 69624
rect 74210 69606 74262 69658
rect 74274 69606 74326 69658
rect 74338 69606 74390 69658
rect 74402 69606 74454 69658
rect 74466 69606 74518 69658
rect 71858 69062 71910 69114
rect 71922 69062 71974 69114
rect 71986 69062 72038 69114
rect 72050 69062 72102 69114
rect 72114 69062 72166 69114
rect 64880 68892 64932 68944
rect 66536 68892 66588 68944
rect 74210 68518 74262 68570
rect 74274 68518 74326 68570
rect 74338 68518 74390 68570
rect 74402 68518 74454 68570
rect 74466 68518 74518 68570
rect 71858 67974 71910 68026
rect 71922 67974 71974 68026
rect 71986 67974 72038 68026
rect 72050 67974 72102 68026
rect 72114 67974 72166 68026
rect 65892 67804 65944 67856
rect 63500 67718 63552 67770
rect 74210 67430 74262 67482
rect 74274 67430 74326 67482
rect 74338 67430 74390 67482
rect 74402 67430 74454 67482
rect 74466 67430 74518 67482
rect 71858 66886 71910 66938
rect 71922 66886 71974 66938
rect 71986 66886 72038 66938
rect 72050 66886 72102 66938
rect 72114 66886 72166 66938
rect 64880 66444 64932 66496
rect 74210 66342 74262 66394
rect 74274 66342 74326 66394
rect 74338 66342 74390 66394
rect 74402 66342 74454 66394
rect 74466 66342 74518 66394
rect 71858 65798 71910 65850
rect 71922 65798 71974 65850
rect 71986 65798 72038 65850
rect 72050 65798 72102 65850
rect 72114 65798 72166 65850
rect 65432 65628 65484 65680
rect 70400 65560 70452 65612
rect 74210 65254 74262 65306
rect 74274 65254 74326 65306
rect 74338 65254 74390 65306
rect 74402 65254 74454 65306
rect 74466 65254 74518 65306
rect 71858 64710 71910 64762
rect 71922 64710 71974 64762
rect 71986 64710 72038 64762
rect 72050 64710 72102 64762
rect 72114 64710 72166 64762
rect 64880 64268 64932 64320
rect 74210 64166 74262 64218
rect 74274 64166 74326 64218
rect 74338 64166 74390 64218
rect 74402 64166 74454 64218
rect 74466 64166 74518 64218
rect 71858 63622 71910 63674
rect 71922 63622 71974 63674
rect 71986 63622 72038 63674
rect 72050 63622 72102 63674
rect 72114 63622 72166 63674
rect 65340 63520 65392 63572
rect 65708 63180 65760 63232
rect 74210 63078 74262 63130
rect 74274 63078 74326 63130
rect 74338 63078 74390 63130
rect 74402 63078 74454 63130
rect 74466 63078 74518 63130
rect 71858 62534 71910 62586
rect 71922 62534 71974 62586
rect 71986 62534 72038 62586
rect 72050 62534 72102 62586
rect 72114 62534 72166 62586
rect 64880 62092 64932 62144
rect 74210 61990 74262 62042
rect 74274 61990 74326 62042
rect 74338 61990 74390 62042
rect 74402 61990 74454 62042
rect 74466 61990 74518 62042
rect 71858 61446 71910 61498
rect 71922 61446 71974 61498
rect 71986 61446 72038 61498
rect 72050 61446 72102 61498
rect 72114 61446 72166 61498
rect 66076 61276 66128 61328
rect 63592 60868 63644 60920
rect 74210 60902 74262 60954
rect 74274 60902 74326 60954
rect 74338 60902 74390 60954
rect 74402 60902 74454 60954
rect 74466 60902 74518 60954
rect 71858 60358 71910 60410
rect 71922 60358 71974 60410
rect 71986 60358 72038 60410
rect 72050 60358 72102 60410
rect 72114 60358 72166 60410
rect 64880 60256 64932 60308
rect 74210 59814 74262 59866
rect 74274 59814 74326 59866
rect 74338 59814 74390 59866
rect 74402 59814 74454 59866
rect 74466 59814 74518 59866
rect 71858 59270 71910 59322
rect 71922 59270 71974 59322
rect 71986 59270 72038 59322
rect 72050 59270 72102 59322
rect 72114 59270 72166 59322
rect 65156 59100 65208 59152
rect 69020 59032 69072 59084
rect 74210 58726 74262 58778
rect 74274 58726 74326 58778
rect 74338 58726 74390 58778
rect 74402 58726 74454 58778
rect 74466 58726 74518 58778
rect 71858 58182 71910 58234
rect 71922 58182 71974 58234
rect 71986 58182 72038 58234
rect 72050 58182 72102 58234
rect 72114 58182 72166 58234
rect 64880 58012 64932 58064
rect 74210 57638 74262 57690
rect 74274 57638 74326 57690
rect 74338 57638 74390 57690
rect 74402 57638 74454 57690
rect 74466 57638 74518 57690
rect 71858 57094 71910 57146
rect 71922 57094 71974 57146
rect 71986 57094 72038 57146
rect 72050 57094 72102 57146
rect 72114 57094 72166 57146
rect 67548 56924 67600 56976
rect 70492 56856 70544 56908
rect 74210 56550 74262 56602
rect 74274 56550 74326 56602
rect 74338 56550 74390 56602
rect 74402 56550 74454 56602
rect 74466 56550 74518 56602
rect 71858 56006 71910 56058
rect 71922 56006 71974 56058
rect 71986 56006 72038 56058
rect 72050 56006 72102 56058
rect 72114 56006 72166 56058
rect 64880 55564 64932 55616
rect 74210 55462 74262 55514
rect 74274 55462 74326 55514
rect 74338 55462 74390 55514
rect 74402 55462 74454 55514
rect 74466 55462 74518 55514
rect 71858 54918 71910 54970
rect 71922 54918 71974 54970
rect 71986 54918 72038 54970
rect 72050 54918 72102 54970
rect 72114 54918 72166 54970
rect 67732 54816 67784 54868
rect 65984 54476 66036 54528
rect 74210 54374 74262 54426
rect 74274 54374 74326 54426
rect 74338 54374 74390 54426
rect 74402 54374 74454 54426
rect 74466 54374 74518 54426
rect 71858 53830 71910 53882
rect 71922 53830 71974 53882
rect 71986 53830 72038 53882
rect 72050 53830 72102 53882
rect 72114 53830 72166 53882
rect 64880 53524 64932 53576
rect 74210 53286 74262 53338
rect 74274 53286 74326 53338
rect 74338 53286 74390 53338
rect 74402 53286 74454 53338
rect 74466 53286 74518 53338
rect 66904 53116 66956 53168
rect 71858 52742 71910 52794
rect 71922 52742 71974 52794
rect 71986 52742 72038 52794
rect 72050 52742 72102 52794
rect 72114 52742 72166 52794
rect 66812 52572 66864 52624
rect 63776 52436 63828 52488
rect 65616 52479 65668 52488
rect 65616 52445 65625 52479
rect 65625 52445 65659 52479
rect 65659 52445 65668 52479
rect 65616 52436 65668 52445
rect 74210 52198 74262 52250
rect 74274 52198 74326 52250
rect 74338 52198 74390 52250
rect 74402 52198 74454 52250
rect 74466 52198 74518 52250
rect 65616 52096 65668 52148
rect 71858 51654 71910 51706
rect 71922 51654 71974 51706
rect 71986 51654 72038 51706
rect 72050 51654 72102 51706
rect 72114 51654 72166 51706
rect 64880 51484 64932 51536
rect 66352 51484 66404 51536
rect 74210 51110 74262 51162
rect 74274 51110 74326 51162
rect 74338 51110 74390 51162
rect 74402 51110 74454 51162
rect 74466 51110 74518 51162
rect 71858 50566 71910 50618
rect 71922 50566 71974 50618
rect 71986 50566 72038 50618
rect 72050 50566 72102 50618
rect 72114 50566 72166 50618
rect 67640 50464 67692 50516
rect 63776 50260 63828 50312
rect 74210 50022 74262 50074
rect 74274 50022 74326 50074
rect 74338 50022 74390 50074
rect 74402 50022 74454 50074
rect 74466 50022 74518 50074
rect 71858 49478 71910 49530
rect 71922 49478 71974 49530
rect 71986 49478 72038 49530
rect 72050 49478 72102 49530
rect 72114 49478 72166 49530
rect 65248 49104 65300 49156
rect 74210 48934 74262 48986
rect 74274 48934 74326 48986
rect 74338 48934 74390 48986
rect 74402 48934 74454 48986
rect 74466 48934 74518 48986
rect 71858 48390 71910 48442
rect 71922 48390 71974 48442
rect 71986 48390 72038 48442
rect 72050 48390 72102 48442
rect 72114 48390 72166 48442
rect 64972 48084 65024 48136
rect 74210 47846 74262 47898
rect 74274 47846 74326 47898
rect 74338 47846 74390 47898
rect 74402 47846 74454 47898
rect 74466 47846 74518 47898
rect 64420 47676 64472 47728
rect 64604 47336 64656 47388
rect 71858 47302 71910 47354
rect 71922 47302 71974 47354
rect 71986 47302 72038 47354
rect 72050 47302 72102 47354
rect 72114 47302 72166 47354
rect 63868 46996 63920 47048
rect 68376 46996 68428 47048
rect 67180 46928 67232 46980
rect 74210 46758 74262 46810
rect 74274 46758 74326 46810
rect 74338 46758 74390 46810
rect 74402 46758 74454 46810
rect 74466 46758 74518 46810
rect 71858 46214 71910 46266
rect 71922 46214 71974 46266
rect 71986 46214 72038 46266
rect 72050 46214 72102 46266
rect 72114 46214 72166 46266
rect 64052 45908 64104 45960
rect 64144 45704 64196 45756
rect 74210 45670 74262 45722
rect 74274 45670 74326 45722
rect 74338 45670 74390 45722
rect 74402 45670 74454 45722
rect 74466 45670 74518 45722
rect 63960 45228 64012 45280
rect 71858 45126 71910 45178
rect 71922 45126 71974 45178
rect 71986 45126 72038 45178
rect 72050 45126 72102 45178
rect 72114 45126 72166 45178
rect 64972 44820 65024 44872
rect 74210 44582 74262 44634
rect 74274 44582 74326 44634
rect 74338 44582 74390 44634
rect 74402 44582 74454 44634
rect 74466 44582 74518 44634
rect 68192 44480 68244 44532
rect 68284 44412 68336 44464
rect 71858 44038 71910 44090
rect 71922 44038 71974 44090
rect 71986 44038 72038 44090
rect 72050 44038 72102 44090
rect 72114 44038 72166 44090
rect 64236 43800 64288 43852
rect 74210 43494 74262 43546
rect 74274 43494 74326 43546
rect 74338 43494 74390 43546
rect 74402 43494 74454 43546
rect 74466 43494 74518 43546
rect 63776 43256 63828 43308
rect 68560 43052 68612 43104
rect 71858 42950 71910 43002
rect 71922 42950 71974 43002
rect 71986 42950 72038 43002
rect 72050 42950 72102 43002
rect 72114 42950 72166 43002
rect 66996 42712 67048 42764
rect 70032 42644 70084 42696
rect 74210 42406 74262 42458
rect 74274 42406 74326 42458
rect 74338 42406 74390 42458
rect 74402 42406 74454 42458
rect 74466 42406 74518 42458
rect 71858 41862 71910 41914
rect 71922 41862 71974 41914
rect 71986 41862 72038 41914
rect 72050 41862 72102 41914
rect 72114 41862 72166 41914
rect 67088 41803 67140 41812
rect 67088 41769 67097 41803
rect 67097 41769 67131 41803
rect 67131 41769 67140 41803
rect 67088 41760 67140 41769
rect 64880 41692 64932 41744
rect 70124 41556 70176 41608
rect 74210 41318 74262 41370
rect 74274 41318 74326 41370
rect 74338 41318 74390 41370
rect 74402 41318 74454 41370
rect 74466 41318 74518 41370
rect 65248 40944 65300 40996
rect 68652 40876 68704 40928
rect 71858 40774 71910 40826
rect 71922 40774 71974 40826
rect 71986 40774 72038 40826
rect 72050 40774 72102 40826
rect 72114 40774 72166 40826
rect 66444 40715 66496 40724
rect 66444 40681 66453 40715
rect 66453 40681 66487 40715
rect 66487 40681 66496 40715
rect 66444 40672 66496 40681
rect 69204 40468 69256 40520
rect 74210 40230 74262 40282
rect 74274 40230 74326 40282
rect 74338 40230 74390 40282
rect 74402 40230 74454 40282
rect 74466 40230 74518 40282
rect 64880 39788 64932 39840
rect 71858 39686 71910 39738
rect 71922 39686 71974 39738
rect 71986 39686 72038 39738
rect 72050 39686 72102 39738
rect 72114 39686 72166 39738
rect 66260 39584 66312 39636
rect 67456 39380 67508 39432
rect 74210 39142 74262 39194
rect 74274 39142 74326 39194
rect 74338 39142 74390 39194
rect 74402 39142 74454 39194
rect 74466 39142 74518 39194
rect 65248 38768 65300 38820
rect 67916 38700 67968 38752
rect 71858 38598 71910 38650
rect 71922 38598 71974 38650
rect 71986 38598 72038 38650
rect 72050 38598 72102 38650
rect 72114 38598 72166 38650
rect 67824 38496 67876 38548
rect 66996 38292 67048 38344
rect 74210 38054 74262 38106
rect 74274 38054 74326 38106
rect 74338 38054 74390 38106
rect 74402 38054 74454 38106
rect 74466 38054 74518 38106
rect 71858 37510 71910 37562
rect 71922 37510 71974 37562
rect 71986 37510 72038 37562
rect 72050 37510 72102 37562
rect 72114 37510 72166 37562
rect 64880 37340 64932 37392
rect 67272 37204 67324 37256
rect 66628 37136 66680 37188
rect 74210 36966 74262 37018
rect 74274 36966 74326 37018
rect 74338 36966 74390 37018
rect 74402 36966 74454 37018
rect 74466 36966 74518 37018
rect 65800 36524 65852 36576
rect 71858 36422 71910 36474
rect 71922 36422 71974 36474
rect 71986 36422 72038 36474
rect 72050 36422 72102 36474
rect 72114 36422 72166 36474
rect 65524 36320 65576 36372
rect 68100 36252 68152 36304
rect 67364 36116 67416 36168
rect 74210 35878 74262 35930
rect 74274 35878 74326 35930
rect 74338 35878 74390 35930
rect 74402 35878 74454 35930
rect 74466 35878 74518 35930
rect 66536 35751 66588 35760
rect 66536 35717 66545 35751
rect 66545 35717 66579 35751
rect 66579 35717 66588 35751
rect 66536 35708 66588 35717
rect 68008 35640 68060 35692
rect 71858 35334 71910 35386
rect 71922 35334 71974 35386
rect 71986 35334 72038 35386
rect 72050 35334 72102 35386
rect 72114 35334 72166 35386
rect 65892 35232 65944 35284
rect 64880 35164 64932 35216
rect 66628 35028 66680 35080
rect 74210 34790 74262 34842
rect 74274 34790 74326 34842
rect 74338 34790 74390 34842
rect 74402 34790 74454 34842
rect 74466 34790 74518 34842
rect 65248 34484 65300 34536
rect 71858 34246 71910 34298
rect 71922 34246 71974 34298
rect 71986 34246 72038 34298
rect 72050 34246 72102 34298
rect 72114 34246 72166 34298
rect 66904 34187 66956 34196
rect 66904 34153 66913 34187
rect 66913 34153 66947 34187
rect 66947 34153 66956 34187
rect 66904 34144 66956 34153
rect 64788 33940 64840 33992
rect 65616 33915 65668 33924
rect 65616 33881 65625 33915
rect 65625 33881 65659 33915
rect 65659 33881 65668 33915
rect 65616 33872 65668 33881
rect 74210 33702 74262 33754
rect 74274 33702 74326 33754
rect 74338 33702 74390 33754
rect 74402 33702 74454 33754
rect 74466 33702 74518 33754
rect 65432 33600 65484 33652
rect 66720 33396 66772 33448
rect 64880 33260 64932 33312
rect 71858 33158 71910 33210
rect 71922 33158 71974 33210
rect 71986 33158 72038 33210
rect 72050 33158 72102 33210
rect 72114 33158 72166 33210
rect 65340 33056 65392 33108
rect 66444 32988 66496 33040
rect 67548 32988 67600 33040
rect 67548 32852 67600 32904
rect 74210 32614 74262 32666
rect 74274 32614 74326 32666
rect 74338 32614 74390 32666
rect 74402 32614 74454 32666
rect 74466 32614 74518 32666
rect 65340 32172 65392 32224
rect 71858 32070 71910 32122
rect 71922 32070 71974 32122
rect 71986 32070 72038 32122
rect 72050 32070 72102 32122
rect 72114 32070 72166 32122
rect 66076 31968 66128 32020
rect 64420 31764 64472 31816
rect 67088 31764 67140 31816
rect 74210 31526 74262 31578
rect 74274 31526 74326 31578
rect 74338 31526 74390 31578
rect 74402 31526 74454 31578
rect 74466 31526 74518 31578
rect 64880 31084 64932 31136
rect 71858 30982 71910 31034
rect 71922 30982 71974 31034
rect 71986 30982 72038 31034
rect 72050 30982 72102 31034
rect 72114 30982 72166 31034
rect 65156 30880 65208 30932
rect 66812 30676 66864 30728
rect 74210 30438 74262 30490
rect 74274 30438 74326 30490
rect 74338 30438 74390 30490
rect 74402 30438 74454 30490
rect 74466 30438 74518 30490
rect 65432 29996 65484 30048
rect 71858 29894 71910 29946
rect 71922 29894 71974 29946
rect 71986 29894 72038 29946
rect 72050 29894 72102 29946
rect 72114 29894 72166 29946
rect 66444 29792 66496 29844
rect 64328 29588 64380 29640
rect 66444 29588 66496 29640
rect 74210 29350 74262 29402
rect 74274 29350 74326 29402
rect 74338 29350 74390 29402
rect 74402 29350 74454 29402
rect 74466 29350 74518 29402
rect 71858 28806 71910 28858
rect 71922 28806 71974 28858
rect 71986 28806 72038 28858
rect 72050 28806 72102 28858
rect 72114 28806 72166 28858
rect 67732 28704 67784 28756
rect 64880 28636 64932 28688
rect 66260 28543 66312 28552
rect 66260 28509 66269 28543
rect 66269 28509 66303 28543
rect 66303 28509 66312 28543
rect 66260 28500 66312 28509
rect 74210 28262 74262 28314
rect 74274 28262 74326 28314
rect 74338 28262 74390 28314
rect 74402 28262 74454 28314
rect 74466 28262 74518 28314
rect 65892 27820 65944 27872
rect 71858 27718 71910 27770
rect 71922 27718 71974 27770
rect 71986 27718 72038 27770
rect 72050 27718 72102 27770
rect 72114 27718 72166 27770
rect 64512 27616 64564 27668
rect 66536 27548 66588 27600
rect 66996 27412 67048 27464
rect 74210 27174 74262 27226
rect 74274 27174 74326 27226
rect 74338 27174 74390 27226
rect 74402 27174 74454 27226
rect 74466 27174 74518 27226
rect 64880 27004 64932 27056
rect 68836 27004 68888 27056
rect 68744 26936 68796 26988
rect 66352 26911 66404 26920
rect 66352 26877 66361 26911
rect 66361 26877 66395 26911
rect 66395 26877 66404 26911
rect 66352 26868 66404 26877
rect 71858 26630 71910 26682
rect 71922 26630 71974 26682
rect 71986 26630 72038 26682
rect 72050 26630 72102 26682
rect 72114 26630 72166 26682
rect 67640 26528 67692 26580
rect 66536 26324 66588 26376
rect 74210 26086 74262 26138
rect 74274 26086 74326 26138
rect 74338 26086 74390 26138
rect 74402 26086 74454 26138
rect 74466 26086 74518 26138
rect 65616 25644 65668 25696
rect 71858 25542 71910 25594
rect 71922 25542 71974 25594
rect 71986 25542 72038 25594
rect 72050 25542 72102 25594
rect 72114 25542 72166 25594
rect 63776 25236 63828 25288
rect 74210 24998 74262 25050
rect 74274 24998 74326 25050
rect 74338 24998 74390 25050
rect 74402 24998 74454 25050
rect 74466 24998 74518 25050
rect 71858 24454 71910 24506
rect 71922 24454 71974 24506
rect 71986 24454 72038 24506
rect 72050 24454 72102 24506
rect 72114 24454 72166 24506
rect 68284 24352 68336 24404
rect 65156 24284 65208 24336
rect 66352 24148 66404 24200
rect 74210 23910 74262 23962
rect 74274 23910 74326 23962
rect 74338 23910 74390 23962
rect 74402 23910 74454 23962
rect 74466 23910 74518 23962
rect 64972 23808 65024 23860
rect 66536 23740 66588 23792
rect 66996 23740 67048 23792
rect 66536 23604 66588 23656
rect 66076 23468 66128 23520
rect 71858 23366 71910 23418
rect 71922 23366 71974 23418
rect 71986 23366 72038 23418
rect 72050 23366 72102 23418
rect 72114 23366 72166 23418
rect 68192 23264 68244 23316
rect 68928 23196 68980 23248
rect 66536 23060 66588 23112
rect 74210 22822 74262 22874
rect 74274 22822 74326 22874
rect 74338 22822 74390 22874
rect 74402 22822 74454 22874
rect 74466 22822 74518 22874
rect 71858 22278 71910 22330
rect 71922 22278 71974 22330
rect 71986 22278 72038 22330
rect 72050 22278 72102 22330
rect 72114 22278 72166 22330
rect 65156 22108 65208 22160
rect 74210 21734 74262 21786
rect 74274 21734 74326 21786
rect 74338 21734 74390 21786
rect 74402 21734 74454 21786
rect 74466 21734 74518 21786
rect 70584 21496 70636 21548
rect 71858 21190 71910 21242
rect 71922 21190 71974 21242
rect 71986 21190 72038 21242
rect 72050 21190 72102 21242
rect 72114 21190 72166 21242
rect 67824 21088 67876 21140
rect 74210 20646 74262 20698
rect 74274 20646 74326 20698
rect 74338 20646 74390 20698
rect 74402 20646 74454 20698
rect 74466 20646 74518 20698
rect 65156 20204 65208 20256
rect 71858 20102 71910 20154
rect 71922 20102 71974 20154
rect 71986 20102 72038 20154
rect 72050 20102 72102 20154
rect 72114 20102 72166 20154
rect 74210 19558 74262 19610
rect 74274 19558 74326 19610
rect 74338 19558 74390 19610
rect 74402 19558 74454 19610
rect 74466 19558 74518 19610
rect 65524 19116 65576 19168
rect 71858 19014 71910 19066
rect 71922 19014 71974 19066
rect 71986 19014 72038 19066
rect 72050 19014 72102 19066
rect 72114 19014 72166 19066
rect 64696 18708 64748 18760
rect 74210 18470 74262 18522
rect 74274 18470 74326 18522
rect 74338 18470 74390 18522
rect 74402 18470 74454 18522
rect 74466 18470 74518 18522
rect 65156 17960 65208 18012
rect 71858 17926 71910 17978
rect 71922 17926 71974 17978
rect 71986 17926 72038 17978
rect 72050 17926 72102 17978
rect 72114 17926 72166 17978
rect 74210 17382 74262 17434
rect 74274 17382 74326 17434
rect 74338 17382 74390 17434
rect 74402 17382 74454 17434
rect 74466 17382 74518 17434
rect 70676 17144 70728 17196
rect 71858 16838 71910 16890
rect 71922 16838 71974 16890
rect 71986 16838 72038 16890
rect 72050 16838 72102 16890
rect 72114 16838 72166 16890
rect 63684 16532 63736 16584
rect 74210 16294 74262 16346
rect 74274 16294 74326 16346
rect 74338 16294 74390 16346
rect 74402 16294 74454 16346
rect 74466 16294 74518 16346
rect 71858 15750 71910 15802
rect 71922 15750 71974 15802
rect 71986 15750 72038 15802
rect 72050 15750 72102 15802
rect 72114 15750 72166 15802
rect 65156 15580 65208 15632
rect 74210 15206 74262 15258
rect 74274 15206 74326 15258
rect 74338 15206 74390 15258
rect 74402 15206 74454 15258
rect 74466 15206 74518 15258
rect 65524 14764 65576 14816
rect 71858 14662 71910 14714
rect 71922 14662 71974 14714
rect 71986 14662 72038 14714
rect 72050 14662 72102 14714
rect 72114 14662 72166 14714
rect 67640 14560 67692 14612
rect 74210 14118 74262 14170
rect 74274 14118 74326 14170
rect 74338 14118 74390 14170
rect 74402 14118 74454 14170
rect 74466 14118 74518 14170
rect 65156 13676 65208 13728
rect 71858 13574 71910 13626
rect 71922 13574 71974 13626
rect 71986 13574 72038 13626
rect 72050 13574 72102 13626
rect 72114 13574 72166 13626
rect 74210 13030 74262 13082
rect 74274 13030 74326 13082
rect 74338 13030 74390 13082
rect 74402 13030 74454 13082
rect 74466 13030 74518 13082
rect 64880 12724 64932 12776
rect 67732 12588 67784 12640
rect 71858 12486 71910 12538
rect 71922 12486 71974 12538
rect 71986 12486 72038 12538
rect 72050 12486 72102 12538
rect 72114 12486 72166 12538
rect 63960 12248 64012 12300
rect 64696 12248 64748 12300
rect 74210 11942 74262 11994
rect 74274 11942 74326 11994
rect 74338 11942 74390 11994
rect 74402 11942 74454 11994
rect 74466 11942 74518 11994
rect 71858 11398 71910 11450
rect 71922 11398 71974 11450
rect 71986 11398 72038 11450
rect 72050 11398 72102 11450
rect 72114 11398 72166 11450
rect 64604 11296 64656 11348
rect 64788 11296 64840 11348
rect 65156 11228 65208 11280
rect 65340 11228 65392 11280
rect 64236 11160 64288 11212
rect 64604 11160 64656 11212
rect 64236 11024 64288 11076
rect 67180 11024 67232 11076
rect 74210 10854 74262 10906
rect 74274 10854 74326 10906
rect 74338 10854 74390 10906
rect 74402 10854 74454 10906
rect 74466 10854 74518 10906
rect 64880 10548 64932 10600
rect 65156 10548 65208 10600
rect 64880 10412 64932 10464
rect 63408 10292 63460 10344
rect 71858 10310 71910 10362
rect 71922 10310 71974 10362
rect 71986 10310 72038 10362
rect 72050 10310 72102 10362
rect 72114 10310 72166 10362
rect 74210 9766 74262 9818
rect 74274 9766 74326 9818
rect 74338 9766 74390 9818
rect 74402 9766 74454 9818
rect 74466 9766 74518 9818
rect 71858 9222 71910 9274
rect 71922 9222 71974 9274
rect 71986 9222 72038 9274
rect 72050 9222 72102 9274
rect 72114 9222 72166 9274
rect 65340 9120 65392 9172
rect 74210 8678 74262 8730
rect 74274 8678 74326 8730
rect 74338 8678 74390 8730
rect 74402 8678 74454 8730
rect 74466 8678 74518 8730
rect 71858 8134 71910 8186
rect 71922 8134 71974 8186
rect 71986 8134 72038 8186
rect 72050 8134 72102 8186
rect 72114 8134 72166 8186
rect 59560 7760 59612 7812
rect 64236 7896 64288 7948
rect 61660 7828 61712 7880
rect 63500 7828 63552 7880
rect 62488 7760 62540 7812
rect 64972 7760 65024 7812
rect 52276 7692 52328 7744
rect 63684 7692 63736 7744
rect 56140 7624 56192 7676
rect 63408 7624 63460 7676
rect 56508 7556 56560 7608
rect 63592 7556 63644 7608
rect 74210 7590 74262 7642
rect 74274 7590 74326 7642
rect 74338 7590 74390 7642
rect 74402 7590 74454 7642
rect 74466 7590 74518 7642
rect 48228 7488 48280 7540
rect 64328 7488 64380 7540
rect 59176 7420 59228 7472
rect 68376 7420 68428 7472
rect 62764 7352 62816 7404
rect 65708 7352 65760 7404
rect 63040 7284 63092 7336
rect 65524 7284 65576 7336
rect 60372 7216 60424 7268
rect 64696 7216 64748 7268
rect 60096 7012 60148 7064
rect 65156 7012 65208 7064
rect 71858 7046 71910 7098
rect 71922 7046 71974 7098
rect 71986 7046 72038 7098
rect 72050 7046 72102 7098
rect 72114 7046 72166 7098
rect 55588 6944 55640 6996
rect 55680 6876 55732 6928
rect 48872 6808 48924 6860
rect 56048 6808 56100 6860
rect 60004 6808 60056 6860
rect 65800 6808 65852 6860
rect 66628 6808 66680 6860
rect 68928 6808 68980 6860
rect 27528 6740 27580 6792
rect 64880 6740 64932 6792
rect 65156 6740 65208 6792
rect 66812 6740 66864 6792
rect 23296 6672 23348 6724
rect 70676 6672 70728 6724
rect 24768 6604 24820 6656
rect 70584 6604 70636 6656
rect 25872 6536 25924 6588
rect 62488 6536 62540 6588
rect 63500 6536 63552 6588
rect 64972 6536 65024 6588
rect 28632 6468 28684 6520
rect 46388 6468 46440 6520
rect 54668 6468 54720 6520
rect 59544 6468 59596 6520
rect 59636 6468 59688 6520
rect 63776 6468 63828 6520
rect 64052 6468 64104 6520
rect 64328 6468 64380 6520
rect 74210 6502 74262 6554
rect 74274 6502 74326 6554
rect 74338 6502 74390 6554
rect 74402 6502 74454 6554
rect 74466 6502 74518 6554
rect 29552 6400 29604 6452
rect 47492 6400 47544 6452
rect 49608 6400 49660 6452
rect 63868 6400 63920 6452
rect 64236 6400 64288 6452
rect 66444 6400 66496 6452
rect 23664 6332 23716 6384
rect 32312 6332 32364 6384
rect 48136 6332 48188 6384
rect 64420 6332 64472 6384
rect 65524 6332 65576 6384
rect 66720 6332 66772 6384
rect 26148 6264 26200 6316
rect 34888 6264 34940 6316
rect 53932 6264 53984 6316
rect 59912 6264 59964 6316
rect 60004 6264 60056 6316
rect 67824 6264 67876 6316
rect 27068 6196 27120 6248
rect 45652 6196 45704 6248
rect 51080 6196 51132 6248
rect 55588 6196 55640 6248
rect 24952 6128 25004 6180
rect 44916 6128 44968 6180
rect 47032 6128 47084 6180
rect 55772 6128 55824 6180
rect 46296 6060 46348 6112
rect 64328 6196 64380 6248
rect 64972 6196 65024 6248
rect 66536 6196 66588 6248
rect 56048 6128 56100 6180
rect 64512 6128 64564 6180
rect 55956 6060 56008 6112
rect 63040 6060 63092 6112
rect 63132 6060 63184 6112
rect 67732 6060 67784 6112
rect 71858 5958 71910 6010
rect 71922 5958 71974 6010
rect 71986 5958 72038 6010
rect 72050 5958 72102 6010
rect 72114 5958 72166 6010
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 33324 5856 33376 5908
rect 33876 5856 33928 5908
rect 48964 5856 49016 5908
rect 49608 5899 49660 5908
rect 49608 5865 49617 5899
rect 49617 5865 49651 5899
rect 49651 5865 49660 5899
rect 49608 5856 49660 5865
rect 55680 5856 55732 5908
rect 55772 5856 55824 5908
rect 59820 5856 59872 5908
rect 59912 5856 59964 5908
rect 63040 5856 63092 5908
rect 63316 5856 63368 5908
rect 65432 5856 65484 5908
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 55956 5788 56008 5840
rect 56232 5788 56284 5840
rect 24584 5720 24636 5772
rect 32220 5720 32272 5772
rect 32588 5720 32640 5772
rect 48872 5763 48924 5772
rect 48872 5729 48881 5763
rect 48881 5729 48915 5763
rect 48915 5729 48924 5763
rect 48872 5720 48924 5729
rect 48964 5763 49016 5772
rect 48964 5729 48973 5763
rect 48973 5729 49007 5763
rect 49007 5729 49016 5763
rect 48964 5720 49016 5729
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 25964 5695 26016 5704
rect 25964 5661 25973 5695
rect 25973 5661 26007 5695
rect 26007 5661 26016 5695
rect 25964 5652 26016 5661
rect 26148 5695 26200 5704
rect 26148 5661 26157 5695
rect 26157 5661 26191 5695
rect 26191 5661 26200 5695
rect 26148 5652 26200 5661
rect 40408 5695 40460 5704
rect 40408 5661 40417 5695
rect 40417 5661 40451 5695
rect 40451 5661 40460 5695
rect 40408 5652 40460 5661
rect 41512 5652 41564 5704
rect 43812 5695 43864 5704
rect 43812 5661 43821 5695
rect 43821 5661 43855 5695
rect 43855 5661 43864 5695
rect 43812 5652 43864 5661
rect 44640 5652 44692 5704
rect 44916 5695 44968 5704
rect 44916 5661 44925 5695
rect 44925 5661 44959 5695
rect 44959 5661 44968 5695
rect 44916 5652 44968 5661
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 46296 5695 46348 5704
rect 46296 5661 46305 5695
rect 46305 5661 46339 5695
rect 46339 5661 46348 5695
rect 46296 5652 46348 5661
rect 46388 5695 46440 5704
rect 46388 5661 46397 5695
rect 46397 5661 46431 5695
rect 46431 5661 46440 5695
rect 46388 5652 46440 5661
rect 47032 5695 47084 5704
rect 47032 5661 47041 5695
rect 47041 5661 47075 5695
rect 47075 5661 47084 5695
rect 47032 5652 47084 5661
rect 47492 5695 47544 5704
rect 47492 5661 47501 5695
rect 47501 5661 47535 5695
rect 47535 5661 47544 5695
rect 47492 5652 47544 5661
rect 54668 5720 54720 5772
rect 61476 5788 61528 5840
rect 56508 5763 56560 5772
rect 56508 5729 56517 5763
rect 56517 5729 56551 5763
rect 56551 5729 56560 5763
rect 56508 5720 56560 5729
rect 57796 5763 57848 5772
rect 57796 5729 57805 5763
rect 57805 5729 57839 5763
rect 57839 5729 57848 5763
rect 57796 5720 57848 5729
rect 58164 5763 58216 5772
rect 58164 5729 58173 5763
rect 58173 5729 58207 5763
rect 58207 5729 58216 5763
rect 58164 5720 58216 5729
rect 58256 5720 58308 5772
rect 59636 5720 59688 5772
rect 59728 5763 59780 5772
rect 59728 5729 59737 5763
rect 59737 5729 59771 5763
rect 59771 5729 59780 5763
rect 59728 5720 59780 5729
rect 59820 5720 59872 5772
rect 63868 5788 63920 5840
rect 61660 5763 61712 5772
rect 61660 5729 61669 5763
rect 61669 5729 61703 5763
rect 61703 5729 61712 5763
rect 61660 5720 61712 5729
rect 62948 5763 63000 5772
rect 62948 5729 62957 5763
rect 62957 5729 62991 5763
rect 62991 5729 63000 5763
rect 62948 5720 63000 5729
rect 63040 5720 63092 5772
rect 67640 5788 67692 5840
rect 64052 5720 64104 5772
rect 64604 5720 64656 5772
rect 65064 5763 65116 5772
rect 65064 5729 65073 5763
rect 65073 5729 65107 5763
rect 65107 5729 65116 5763
rect 65064 5720 65116 5729
rect 66168 5763 66220 5772
rect 66168 5729 66177 5763
rect 66177 5729 66211 5763
rect 66211 5729 66220 5763
rect 66168 5720 66220 5729
rect 68468 5763 68520 5772
rect 68468 5729 68477 5763
rect 68477 5729 68511 5763
rect 68511 5729 68520 5763
rect 68468 5720 68520 5729
rect 37004 5627 37056 5636
rect 37004 5593 37013 5627
rect 37013 5593 37047 5627
rect 37047 5593 37056 5627
rect 37004 5584 37056 5593
rect 47860 5584 47912 5636
rect 31668 5516 31720 5568
rect 35900 5516 35952 5568
rect 41696 5559 41748 5568
rect 41696 5525 41705 5559
rect 41705 5525 41739 5559
rect 41739 5525 41748 5559
rect 41696 5516 41748 5525
rect 50436 5695 50488 5704
rect 50436 5661 50445 5695
rect 50445 5661 50479 5695
rect 50479 5661 50488 5695
rect 50436 5652 50488 5661
rect 51264 5695 51316 5704
rect 51264 5661 51273 5695
rect 51273 5661 51307 5695
rect 51307 5661 51316 5695
rect 51264 5652 51316 5661
rect 52276 5652 52328 5704
rect 52644 5695 52696 5704
rect 52644 5661 52653 5695
rect 52653 5661 52687 5695
rect 52687 5661 52696 5695
rect 52644 5652 52696 5661
rect 53380 5695 53432 5704
rect 53380 5661 53389 5695
rect 53389 5661 53423 5695
rect 53423 5661 53432 5695
rect 53380 5652 53432 5661
rect 53932 5652 53984 5704
rect 54576 5652 54628 5704
rect 55312 5695 55364 5704
rect 55312 5661 55321 5695
rect 55321 5661 55355 5695
rect 55355 5661 55364 5695
rect 55312 5652 55364 5661
rect 56140 5652 56192 5704
rect 56324 5695 56376 5704
rect 56324 5661 56333 5695
rect 56333 5661 56367 5695
rect 56367 5661 56376 5695
rect 56324 5652 56376 5661
rect 61108 5652 61160 5704
rect 48044 5584 48096 5636
rect 61016 5584 61068 5636
rect 48136 5559 48188 5568
rect 48136 5525 48145 5559
rect 48145 5525 48179 5559
rect 48179 5525 48188 5559
rect 48136 5516 48188 5525
rect 58256 5516 58308 5568
rect 59452 5516 59504 5568
rect 59544 5516 59596 5568
rect 64052 5584 64104 5636
rect 61200 5516 61252 5568
rect 61476 5516 61528 5568
rect 63132 5516 63184 5568
rect 63224 5516 63276 5568
rect 63408 5516 63460 5568
rect 68836 5584 68888 5636
rect 64788 5516 64840 5568
rect 66444 5516 66496 5568
rect 68100 5559 68152 5568
rect 68100 5525 68109 5559
rect 68109 5525 68143 5559
rect 68143 5525 68152 5559
rect 68100 5516 68152 5525
rect 4210 5414 4262 5466
rect 4274 5414 4326 5466
rect 4338 5414 4390 5466
rect 4402 5414 4454 5466
rect 4466 5414 4518 5466
rect 14210 5414 14262 5466
rect 14274 5414 14326 5466
rect 14338 5414 14390 5466
rect 14402 5414 14454 5466
rect 14466 5414 14518 5466
rect 24210 5414 24262 5466
rect 24274 5414 24326 5466
rect 24338 5414 24390 5466
rect 24402 5414 24454 5466
rect 24466 5414 24518 5466
rect 34210 5414 34262 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 44210 5414 44262 5466
rect 44274 5414 44326 5466
rect 44338 5414 44390 5466
rect 44402 5414 44454 5466
rect 44466 5414 44518 5466
rect 54210 5414 54262 5466
rect 54274 5414 54326 5466
rect 54338 5414 54390 5466
rect 54402 5414 54454 5466
rect 54466 5414 54518 5466
rect 64210 5414 64262 5466
rect 64274 5414 64326 5466
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 74210 5414 74262 5466
rect 74274 5414 74326 5466
rect 74338 5414 74390 5466
rect 74402 5414 74454 5466
rect 74466 5414 74518 5466
rect 23940 5176 23992 5228
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 24584 5108 24636 5160
rect 25412 5151 25464 5160
rect 25412 5117 25421 5151
rect 25421 5117 25455 5151
rect 25455 5117 25464 5151
rect 25412 5108 25464 5117
rect 25964 5312 26016 5364
rect 27804 5312 27856 5364
rect 36820 5312 36872 5364
rect 41052 5355 41104 5364
rect 41052 5321 41061 5355
rect 41061 5321 41095 5355
rect 41095 5321 41104 5355
rect 41052 5312 41104 5321
rect 41144 5312 41196 5364
rect 54760 5312 54812 5364
rect 27620 5244 27672 5296
rect 27436 5176 27488 5228
rect 23480 5040 23532 5092
rect 25780 5083 25832 5092
rect 25780 5049 25789 5083
rect 25789 5049 25823 5083
rect 25823 5049 25832 5083
rect 25780 5040 25832 5049
rect 26332 5151 26384 5160
rect 26332 5117 26341 5151
rect 26341 5117 26375 5151
rect 26375 5117 26384 5151
rect 26332 5108 26384 5117
rect 27160 5108 27212 5160
rect 27528 5151 27580 5160
rect 27528 5117 27537 5151
rect 27537 5117 27571 5151
rect 27571 5117 27580 5151
rect 27528 5108 27580 5117
rect 27804 5176 27856 5228
rect 28080 5244 28132 5296
rect 31208 5244 31260 5296
rect 27252 5040 27304 5092
rect 28264 5040 28316 5092
rect 28448 5151 28500 5160
rect 28448 5117 28457 5151
rect 28457 5117 28491 5151
rect 28491 5117 28500 5151
rect 28448 5108 28500 5117
rect 29092 5151 29144 5160
rect 29092 5117 29101 5151
rect 29101 5117 29135 5151
rect 29135 5117 29144 5151
rect 29092 5108 29144 5117
rect 29736 5151 29788 5160
rect 29736 5117 29745 5151
rect 29745 5117 29779 5151
rect 29779 5117 29788 5151
rect 29736 5108 29788 5117
rect 30288 5219 30340 5228
rect 30288 5185 30297 5219
rect 30297 5185 30331 5219
rect 30331 5185 30340 5219
rect 30288 5176 30340 5185
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 31392 5176 31444 5228
rect 40960 5176 41012 5228
rect 54668 5244 54720 5296
rect 41696 5176 41748 5228
rect 40408 5151 40460 5160
rect 40408 5117 40417 5151
rect 40417 5117 40451 5151
rect 40451 5117 40460 5151
rect 40408 5108 40460 5117
rect 40592 5040 40644 5092
rect 42708 5108 42760 5160
rect 44640 5040 44692 5092
rect 26148 4972 26200 5024
rect 26240 5015 26292 5024
rect 26240 4981 26249 5015
rect 26249 4981 26283 5015
rect 26283 4981 26292 5015
rect 26240 4972 26292 4981
rect 26700 5015 26752 5024
rect 26700 4981 26709 5015
rect 26709 4981 26743 5015
rect 26743 4981 26752 5015
rect 26700 4972 26752 4981
rect 28540 4972 28592 5024
rect 28724 5015 28776 5024
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 29368 5015 29420 5024
rect 29368 4981 29377 5015
rect 29377 4981 29411 5015
rect 29411 4981 29420 5015
rect 29368 4972 29420 4981
rect 29460 4972 29512 5024
rect 30472 5015 30524 5024
rect 30472 4981 30481 5015
rect 30481 4981 30515 5015
rect 30515 4981 30524 5015
rect 30472 4972 30524 4981
rect 33048 4972 33100 5024
rect 46204 5219 46256 5228
rect 46204 5185 46213 5219
rect 46213 5185 46247 5219
rect 46247 5185 46256 5219
rect 46204 5176 46256 5185
rect 46296 5219 46348 5228
rect 46296 5185 46305 5219
rect 46305 5185 46339 5219
rect 46339 5185 46348 5219
rect 46296 5176 46348 5185
rect 46572 5151 46624 5160
rect 46572 5117 46581 5151
rect 46581 5117 46615 5151
rect 46615 5117 46624 5151
rect 46572 5108 46624 5117
rect 53012 5176 53064 5228
rect 60648 5312 60700 5364
rect 55036 5244 55088 5296
rect 65892 5312 65944 5364
rect 47216 5040 47268 5092
rect 46020 5015 46072 5024
rect 46020 4981 46029 5015
rect 46029 4981 46063 5015
rect 46063 4981 46072 5015
rect 46020 4972 46072 4981
rect 47124 4972 47176 5024
rect 47492 5151 47544 5160
rect 47492 5117 47501 5151
rect 47501 5117 47535 5151
rect 47535 5117 47544 5151
rect 47492 5108 47544 5117
rect 48228 5108 48280 5160
rect 49148 5151 49200 5160
rect 49148 5117 49157 5151
rect 49157 5117 49191 5151
rect 49191 5117 49200 5151
rect 49148 5108 49200 5117
rect 50988 5108 51040 5160
rect 53288 5151 53340 5160
rect 53288 5117 53297 5151
rect 53297 5117 53331 5151
rect 53331 5117 53340 5151
rect 53288 5108 53340 5117
rect 56324 5176 56376 5228
rect 56416 5176 56468 5228
rect 65340 5244 65392 5296
rect 69664 5244 69716 5296
rect 61292 5176 61344 5228
rect 55128 5108 55180 5160
rect 65616 5108 65668 5160
rect 69940 5108 69992 5160
rect 47400 5040 47452 5092
rect 49516 4972 49568 5024
rect 52920 5015 52972 5024
rect 52920 4981 52929 5015
rect 52929 4981 52963 5015
rect 52963 4981 52972 5015
rect 52920 4972 52972 4981
rect 54668 4972 54720 5024
rect 55956 5040 56008 5092
rect 66076 5040 66128 5092
rect 69756 5040 69808 5092
rect 68192 4972 68244 5024
rect 69848 4972 69900 5024
rect 71412 4972 71464 5024
rect 73252 5015 73304 5024
rect 73252 4981 73261 5015
rect 73261 4981 73295 5015
rect 73295 4981 73304 5015
rect 73252 4972 73304 4981
rect 1858 4870 1910 4922
rect 1922 4870 1974 4922
rect 1986 4870 2038 4922
rect 2050 4870 2102 4922
rect 2114 4870 2166 4922
rect 11858 4870 11910 4922
rect 11922 4870 11974 4922
rect 11986 4870 12038 4922
rect 12050 4870 12102 4922
rect 12114 4870 12166 4922
rect 21858 4870 21910 4922
rect 21922 4870 21974 4922
rect 21986 4870 22038 4922
rect 22050 4870 22102 4922
rect 22114 4870 22166 4922
rect 31858 4870 31910 4922
rect 31922 4870 31974 4922
rect 31986 4870 32038 4922
rect 32050 4870 32102 4922
rect 32114 4870 32166 4922
rect 41858 4870 41910 4922
rect 41922 4870 41974 4922
rect 41986 4870 42038 4922
rect 42050 4870 42102 4922
rect 42114 4870 42166 4922
rect 51858 4870 51910 4922
rect 51922 4870 51974 4922
rect 51986 4870 52038 4922
rect 52050 4870 52102 4922
rect 52114 4870 52166 4922
rect 61858 4870 61910 4922
rect 61922 4870 61974 4922
rect 61986 4870 62038 4922
rect 62050 4870 62102 4922
rect 62114 4870 62166 4922
rect 71858 4870 71910 4922
rect 71922 4870 71974 4922
rect 71986 4870 72038 4922
rect 72050 4870 72102 4922
rect 72114 4870 72166 4922
rect 26240 4768 26292 4820
rect 30012 4768 30064 4820
rect 31024 4768 31076 4820
rect 40592 4768 40644 4820
rect 25412 4700 25464 4752
rect 24584 4632 24636 4684
rect 31392 4632 31444 4684
rect 35072 4700 35124 4752
rect 41696 4700 41748 4752
rect 43352 4632 43404 4684
rect 44732 4768 44784 4820
rect 46020 4768 46072 4820
rect 60096 4768 60148 4820
rect 61108 4811 61160 4820
rect 61108 4777 61117 4811
rect 61117 4777 61151 4811
rect 61151 4777 61160 4811
rect 61108 4768 61160 4777
rect 45100 4700 45152 4752
rect 44732 4632 44784 4684
rect 48964 4632 49016 4684
rect 27620 4564 27672 4616
rect 33784 4564 33836 4616
rect 33968 4607 34020 4616
rect 33968 4573 33977 4607
rect 33977 4573 34011 4607
rect 34011 4573 34020 4607
rect 33968 4564 34020 4573
rect 34060 4564 34112 4616
rect 41236 4607 41288 4616
rect 41236 4573 41245 4607
rect 41245 4573 41279 4607
rect 41279 4573 41288 4607
rect 41236 4564 41288 4573
rect 41696 4564 41748 4616
rect 43536 4564 43588 4616
rect 26700 4496 26752 4548
rect 29276 4496 29328 4548
rect 29736 4496 29788 4548
rect 34704 4496 34756 4548
rect 46296 4564 46348 4616
rect 46664 4564 46716 4616
rect 46756 4607 46808 4616
rect 46756 4573 46765 4607
rect 46765 4573 46799 4607
rect 46799 4573 46808 4607
rect 46756 4564 46808 4573
rect 46848 4607 46900 4616
rect 46848 4573 46857 4607
rect 46857 4573 46891 4607
rect 46891 4573 46900 4607
rect 46848 4564 46900 4573
rect 46940 4496 46992 4548
rect 53012 4700 53064 4752
rect 60372 4700 60424 4752
rect 62672 4700 62724 4752
rect 49424 4564 49476 4616
rect 61384 4632 61436 4684
rect 69020 4632 69072 4684
rect 61292 4564 61344 4616
rect 62672 4564 62724 4616
rect 67916 4564 67968 4616
rect 26148 4428 26200 4480
rect 29644 4428 29696 4480
rect 33784 4428 33836 4480
rect 34796 4428 34848 4480
rect 35716 4428 35768 4480
rect 42524 4428 42576 4480
rect 42616 4471 42668 4480
rect 42616 4437 42625 4471
rect 42625 4437 42659 4471
rect 42659 4437 42668 4471
rect 42616 4428 42668 4437
rect 43996 4471 44048 4480
rect 43996 4437 44005 4471
rect 44005 4437 44039 4471
rect 44039 4437 44048 4471
rect 43996 4428 44048 4437
rect 45928 4428 45980 4480
rect 49056 4428 49108 4480
rect 60740 4496 60792 4548
rect 62764 4496 62816 4548
rect 68652 4496 68704 4548
rect 60832 4428 60884 4480
rect 61016 4428 61068 4480
rect 68560 4428 68612 4480
rect 4210 4326 4262 4378
rect 4274 4326 4326 4378
rect 4338 4326 4390 4378
rect 4402 4326 4454 4378
rect 4466 4326 4518 4378
rect 14210 4326 14262 4378
rect 14274 4326 14326 4378
rect 14338 4326 14390 4378
rect 14402 4326 14454 4378
rect 14466 4326 14518 4378
rect 24210 4326 24262 4378
rect 24274 4326 24326 4378
rect 24338 4326 24390 4378
rect 24402 4326 24454 4378
rect 24466 4326 24518 4378
rect 34210 4326 34262 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 44210 4326 44262 4378
rect 44274 4326 44326 4378
rect 44338 4326 44390 4378
rect 44402 4326 44454 4378
rect 44466 4326 44518 4378
rect 54210 4326 54262 4378
rect 54274 4326 54326 4378
rect 54338 4326 54390 4378
rect 54402 4326 54454 4378
rect 54466 4326 54518 4378
rect 64210 4326 64262 4378
rect 64274 4326 64326 4378
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 74210 4326 74262 4378
rect 74274 4326 74326 4378
rect 74338 4326 74390 4378
rect 74402 4326 74454 4378
rect 74466 4326 74518 4378
rect 26332 4224 26384 4276
rect 63500 4224 63552 4276
rect 19064 4088 19116 4140
rect 20260 4088 20312 4140
rect 27620 4131 27672 4140
rect 27620 4097 27629 4131
rect 27629 4097 27663 4131
rect 27663 4097 27672 4131
rect 27620 4088 27672 4097
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 31392 4088 31444 4140
rect 33048 4156 33100 4208
rect 33784 4088 33836 4140
rect 34704 4131 34756 4140
rect 34704 4097 34713 4131
rect 34713 4097 34747 4131
rect 34747 4097 34756 4131
rect 34704 4088 34756 4097
rect 34796 4088 34848 4140
rect 43996 4156 44048 4208
rect 49424 4156 49476 4208
rect 49516 4156 49568 4208
rect 53288 4156 53340 4208
rect 70492 4156 70544 4208
rect 41696 4020 41748 4072
rect 42616 4020 42668 4072
rect 46940 4020 46992 4072
rect 56416 4088 56468 4140
rect 61108 4088 61160 4140
rect 67548 4088 67600 4140
rect 64972 4020 65024 4072
rect 17868 3952 17920 4004
rect 40408 3952 40460 4004
rect 42524 3952 42576 4004
rect 45100 3952 45152 4004
rect 54024 3952 54076 4004
rect 54576 3952 54628 4004
rect 60832 3952 60884 4004
rect 62764 3952 62816 4004
rect 23572 3884 23624 3936
rect 27620 3884 27672 3936
rect 27712 3927 27764 3936
rect 27712 3893 27721 3927
rect 27721 3893 27755 3927
rect 27755 3893 27764 3927
rect 27712 3884 27764 3893
rect 33968 3884 34020 3936
rect 35992 3884 36044 3936
rect 49148 3884 49200 3936
rect 1858 3782 1910 3834
rect 1922 3782 1974 3834
rect 1986 3782 2038 3834
rect 2050 3782 2102 3834
rect 2114 3782 2166 3834
rect 11858 3782 11910 3834
rect 11922 3782 11974 3834
rect 11986 3782 12038 3834
rect 12050 3782 12102 3834
rect 12114 3782 12166 3834
rect 21858 3782 21910 3834
rect 21922 3782 21974 3834
rect 21986 3782 22038 3834
rect 22050 3782 22102 3834
rect 22114 3782 22166 3834
rect 31858 3782 31910 3834
rect 31922 3782 31974 3834
rect 31986 3782 32038 3834
rect 32050 3782 32102 3834
rect 32114 3782 32166 3834
rect 41858 3782 41910 3834
rect 41922 3782 41974 3834
rect 41986 3782 42038 3834
rect 42050 3782 42102 3834
rect 42114 3782 42166 3834
rect 51858 3782 51910 3834
rect 51922 3782 51974 3834
rect 51986 3782 52038 3834
rect 52050 3782 52102 3834
rect 52114 3782 52166 3834
rect 61858 3782 61910 3834
rect 61922 3782 61974 3834
rect 61986 3782 62038 3834
rect 62050 3782 62102 3834
rect 62114 3782 62166 3834
rect 71858 3782 71910 3834
rect 71922 3782 71974 3834
rect 71986 3782 72038 3834
rect 72050 3782 72102 3834
rect 72114 3782 72166 3834
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 26056 3723 26108 3732
rect 26056 3689 26065 3723
rect 26065 3689 26099 3723
rect 26099 3689 26108 3723
rect 26056 3680 26108 3689
rect 29736 3680 29788 3732
rect 31300 3680 31352 3732
rect 32404 3723 32456 3732
rect 32404 3689 32413 3723
rect 32413 3689 32447 3723
rect 32447 3689 32456 3723
rect 32404 3680 32456 3689
rect 20628 3544 20680 3596
rect 24952 3587 25004 3596
rect 24952 3553 24961 3587
rect 24961 3553 24995 3587
rect 24995 3553 25004 3587
rect 24952 3544 25004 3553
rect 33416 3680 33468 3732
rect 47492 3680 47544 3732
rect 58532 3680 58584 3732
rect 61292 3680 61344 3732
rect 41236 3612 41288 3664
rect 42248 3612 42300 3664
rect 52644 3612 52696 3664
rect 55772 3612 55824 3664
rect 66260 3612 66312 3664
rect 28816 3544 28868 3596
rect 18236 3476 18288 3528
rect 20536 3476 20588 3528
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 22468 3476 22520 3528
rect 23572 3476 23624 3528
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 25780 3519 25832 3528
rect 25780 3485 25789 3519
rect 25789 3485 25823 3519
rect 25823 3485 25832 3519
rect 25780 3476 25832 3485
rect 23112 3340 23164 3392
rect 23296 3383 23348 3392
rect 23296 3349 23305 3383
rect 23305 3349 23339 3383
rect 23339 3349 23348 3383
rect 23296 3340 23348 3349
rect 25872 3451 25924 3460
rect 25872 3417 25881 3451
rect 25881 3417 25915 3451
rect 25915 3417 25924 3451
rect 25872 3408 25924 3417
rect 27988 3476 28040 3528
rect 28724 3476 28776 3528
rect 31392 3544 31444 3596
rect 26148 3408 26200 3460
rect 27712 3451 27764 3460
rect 27712 3417 27721 3451
rect 27721 3417 27755 3451
rect 27755 3417 27764 3451
rect 27712 3408 27764 3417
rect 28172 3408 28224 3460
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 29000 3408 29052 3460
rect 31668 3519 31720 3528
rect 31668 3485 31677 3519
rect 31677 3485 31711 3519
rect 31711 3485 31720 3519
rect 31668 3476 31720 3485
rect 32404 3544 32456 3596
rect 39764 3544 39816 3596
rect 51540 3544 51592 3596
rect 66352 3544 66404 3596
rect 32220 3519 32272 3528
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 32312 3476 32364 3528
rect 33048 3476 33100 3528
rect 38016 3476 38068 3528
rect 44824 3476 44876 3528
rect 58532 3476 58584 3528
rect 60740 3476 60792 3528
rect 67088 3476 67140 3528
rect 44640 3408 44692 3460
rect 48228 3408 48280 3460
rect 66996 3408 67048 3460
rect 27804 3340 27856 3392
rect 27896 3383 27948 3392
rect 27896 3349 27905 3383
rect 27905 3349 27939 3383
rect 27939 3349 27948 3383
rect 27896 3340 27948 3349
rect 27988 3340 28040 3392
rect 31024 3340 31076 3392
rect 32680 3340 32732 3392
rect 36912 3340 36964 3392
rect 37004 3340 37056 3392
rect 47492 3340 47544 3392
rect 4210 3238 4262 3290
rect 4274 3238 4326 3290
rect 4338 3238 4390 3290
rect 4402 3238 4454 3290
rect 4466 3238 4518 3290
rect 14210 3238 14262 3290
rect 14274 3238 14326 3290
rect 14338 3238 14390 3290
rect 14402 3238 14454 3290
rect 14466 3238 14518 3290
rect 24210 3238 24262 3290
rect 24274 3238 24326 3290
rect 24338 3238 24390 3290
rect 24402 3238 24454 3290
rect 24466 3238 24518 3290
rect 34210 3238 34262 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 44210 3238 44262 3290
rect 44274 3238 44326 3290
rect 44338 3238 44390 3290
rect 44402 3238 44454 3290
rect 44466 3238 44518 3290
rect 54210 3238 54262 3290
rect 54274 3238 54326 3290
rect 54338 3238 54390 3290
rect 54402 3238 54454 3290
rect 54466 3238 54518 3290
rect 64210 3238 64262 3290
rect 64274 3238 64326 3290
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 74210 3238 74262 3290
rect 74274 3238 74326 3290
rect 74338 3238 74390 3290
rect 74402 3238 74454 3290
rect 74466 3238 74518 3290
rect 20536 3179 20588 3188
rect 20536 3145 20545 3179
rect 20545 3145 20579 3179
rect 20579 3145 20588 3179
rect 20536 3136 20588 3145
rect 20904 3179 20956 3188
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 24860 3136 24912 3188
rect 25780 3136 25832 3188
rect 27712 3136 27764 3188
rect 29552 3136 29604 3188
rect 17868 3111 17920 3120
rect 17868 3077 17877 3111
rect 17877 3077 17911 3111
rect 17911 3077 17920 3111
rect 17868 3068 17920 3077
rect 22836 3068 22888 3120
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 19340 3000 19392 3052
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 20720 3000 20772 3052
rect 18696 2932 18748 2984
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 20628 2864 20680 2916
rect 21732 2975 21784 2984
rect 21732 2941 21741 2975
rect 21741 2941 21775 2975
rect 21775 2941 21784 2975
rect 21732 2932 21784 2941
rect 26056 3068 26108 3120
rect 23112 3043 23164 3052
rect 23112 3009 23121 3043
rect 23121 3009 23155 3043
rect 23155 3009 23164 3043
rect 23112 3000 23164 3009
rect 29368 3068 29420 3120
rect 33416 3136 33468 3188
rect 33232 3068 33284 3120
rect 23020 2932 23072 2984
rect 24032 2932 24084 2984
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 22284 2864 22336 2916
rect 22836 2864 22888 2916
rect 26148 2864 26200 2916
rect 26976 3000 27028 3052
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 28908 3000 28960 3052
rect 27068 2975 27120 2984
rect 27068 2941 27077 2975
rect 27077 2941 27111 2975
rect 27111 2941 27120 2975
rect 27068 2932 27120 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 28724 2932 28776 2984
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 29552 3043 29604 3052
rect 29552 3009 29561 3043
rect 29561 3009 29595 3043
rect 29595 3009 29604 3043
rect 29552 3000 29604 3009
rect 29644 3000 29696 3052
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 32312 3000 32364 3052
rect 32588 3043 32640 3052
rect 32588 3009 32597 3043
rect 32597 3009 32631 3043
rect 32631 3009 32640 3043
rect 32588 3000 32640 3009
rect 33140 3000 33192 3052
rect 33324 3043 33376 3052
rect 33324 3009 33333 3043
rect 33333 3009 33367 3043
rect 33367 3009 33376 3043
rect 33324 3000 33376 3009
rect 29460 2864 29512 2916
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 22560 2796 22612 2848
rect 24952 2839 25004 2848
rect 24952 2805 24961 2839
rect 24961 2805 24995 2839
rect 24995 2805 25004 2839
rect 24952 2796 25004 2805
rect 25964 2839 26016 2848
rect 25964 2805 25973 2839
rect 25973 2805 26007 2839
rect 26007 2805 26016 2839
rect 25964 2796 26016 2805
rect 26516 2839 26568 2848
rect 26516 2805 26525 2839
rect 26525 2805 26559 2839
rect 26559 2805 26568 2839
rect 26516 2796 26568 2805
rect 28080 2796 28132 2848
rect 30196 2932 30248 2984
rect 30932 2975 30984 2984
rect 30932 2941 30941 2975
rect 30941 2941 30975 2975
rect 30975 2941 30984 2975
rect 30932 2932 30984 2941
rect 32220 2975 32272 2984
rect 32220 2941 32229 2975
rect 32229 2941 32263 2975
rect 32263 2941 32272 2975
rect 32220 2932 32272 2941
rect 34796 3068 34848 3120
rect 33784 3043 33836 3052
rect 33784 3009 33793 3043
rect 33793 3009 33827 3043
rect 33827 3009 33836 3043
rect 33784 3000 33836 3009
rect 34060 3043 34112 3052
rect 34060 3009 34069 3043
rect 34069 3009 34103 3043
rect 34103 3009 34112 3043
rect 34060 3000 34112 3009
rect 34612 3000 34664 3052
rect 34888 3043 34940 3052
rect 34888 3009 34897 3043
rect 34897 3009 34931 3043
rect 34931 3009 34940 3043
rect 34888 3000 34940 3009
rect 37004 3179 37056 3188
rect 37004 3145 37013 3179
rect 37013 3145 37047 3179
rect 37047 3145 37056 3179
rect 37004 3136 37056 3145
rect 35992 3068 36044 3120
rect 47032 3068 47084 3120
rect 51264 3068 51316 3120
rect 63960 3068 64012 3120
rect 35716 3043 35768 3052
rect 35716 3009 35725 3043
rect 35725 3009 35759 3043
rect 35759 3009 35768 3043
rect 35716 3000 35768 3009
rect 36728 3000 36780 3052
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 36912 3000 36964 3052
rect 42432 3000 42484 3052
rect 45928 3043 45980 3052
rect 45928 3009 45937 3043
rect 45937 3009 45971 3043
rect 45971 3009 45980 3043
rect 45928 3000 45980 3009
rect 47124 3000 47176 3052
rect 49056 3043 49108 3052
rect 49056 3009 49065 3043
rect 49065 3009 49099 3043
rect 49099 3009 49108 3043
rect 49056 3000 49108 3009
rect 52920 3043 52972 3052
rect 52920 3009 52929 3043
rect 52929 3009 52963 3043
rect 52963 3009 52972 3043
rect 52920 3000 52972 3009
rect 53932 3000 53984 3052
rect 54668 3043 54720 3052
rect 54668 3009 54677 3043
rect 54677 3009 54711 3043
rect 54711 3009 54720 3043
rect 54668 3000 54720 3009
rect 56232 3043 56284 3052
rect 56232 3009 56241 3043
rect 56241 3009 56275 3043
rect 56275 3009 56284 3043
rect 56232 3000 56284 3009
rect 57796 3043 57848 3052
rect 57796 3009 57805 3043
rect 57805 3009 57839 3043
rect 57839 3009 57848 3043
rect 57796 3000 57848 3009
rect 59452 3043 59504 3052
rect 59452 3009 59461 3043
rect 59461 3009 59495 3043
rect 59495 3009 59504 3043
rect 59452 3000 59504 3009
rect 61200 3043 61252 3052
rect 61200 3009 61209 3043
rect 61209 3009 61243 3043
rect 61243 3009 61252 3043
rect 61200 3000 61252 3009
rect 63224 3043 63276 3052
rect 63224 3009 63233 3043
rect 63233 3009 63267 3043
rect 63267 3009 63276 3043
rect 63224 3000 63276 3009
rect 64788 3043 64840 3052
rect 64788 3009 64797 3043
rect 64797 3009 64831 3043
rect 64831 3009 64840 3043
rect 64788 3000 64840 3009
rect 66444 3043 66496 3052
rect 66444 3009 66453 3043
rect 66453 3009 66487 3043
rect 66487 3009 66496 3043
rect 66444 3000 66496 3009
rect 68100 3043 68152 3052
rect 68100 3009 68109 3043
rect 68109 3009 68143 3043
rect 68143 3009 68152 3043
rect 68100 3000 68152 3009
rect 69848 3043 69900 3052
rect 69848 3009 69857 3043
rect 69857 3009 69891 3043
rect 69891 3009 69900 3043
rect 69848 3000 69900 3009
rect 71412 3043 71464 3052
rect 71412 3009 71421 3043
rect 71421 3009 71455 3043
rect 71455 3009 71464 3043
rect 71412 3000 71464 3009
rect 73252 3000 73304 3052
rect 42984 2932 43036 2984
rect 33876 2796 33928 2848
rect 35716 2864 35768 2916
rect 44824 2864 44876 2916
rect 50068 2864 50120 2916
rect 44916 2796 44968 2848
rect 47584 2796 47636 2848
rect 52644 2796 52696 2848
rect 53104 2839 53156 2848
rect 53104 2805 53113 2839
rect 53113 2805 53147 2839
rect 53147 2805 53156 2839
rect 53104 2796 53156 2805
rect 55220 2796 55272 2848
rect 56416 2839 56468 2848
rect 56416 2805 56425 2839
rect 56425 2805 56459 2839
rect 56459 2805 56468 2839
rect 56416 2796 56468 2805
rect 57980 2839 58032 2848
rect 57980 2805 57989 2839
rect 57989 2805 58023 2839
rect 58023 2805 58032 2839
rect 57980 2796 58032 2805
rect 60372 2796 60424 2848
rect 61384 2839 61436 2848
rect 61384 2805 61393 2839
rect 61393 2805 61427 2839
rect 61427 2805 61436 2839
rect 61384 2796 61436 2805
rect 63040 2839 63092 2848
rect 63040 2805 63049 2839
rect 63049 2805 63083 2839
rect 63083 2805 63092 2839
rect 63040 2796 63092 2805
rect 64604 2839 64656 2848
rect 64604 2805 64613 2839
rect 64613 2805 64647 2839
rect 64647 2805 64656 2839
rect 64604 2796 64656 2805
rect 66260 2839 66312 2848
rect 66260 2805 66269 2839
rect 66269 2805 66303 2839
rect 66303 2805 66312 2839
rect 66260 2796 66312 2805
rect 68284 2839 68336 2848
rect 68284 2805 68293 2839
rect 68293 2805 68327 2839
rect 68327 2805 68336 2839
rect 68284 2796 68336 2805
rect 69664 2839 69716 2848
rect 69664 2805 69673 2839
rect 69673 2805 69707 2839
rect 69707 2805 69716 2839
rect 69664 2796 69716 2805
rect 71228 2839 71280 2848
rect 71228 2805 71237 2839
rect 71237 2805 71271 2839
rect 71271 2805 71280 2839
rect 71228 2796 71280 2805
rect 73252 2796 73304 2848
rect 1858 2694 1910 2746
rect 1922 2694 1974 2746
rect 1986 2694 2038 2746
rect 2050 2694 2102 2746
rect 2114 2694 2166 2746
rect 11858 2694 11910 2746
rect 11922 2694 11974 2746
rect 11986 2694 12038 2746
rect 12050 2694 12102 2746
rect 12114 2694 12166 2746
rect 21858 2694 21910 2746
rect 21922 2694 21974 2746
rect 21986 2694 22038 2746
rect 22050 2694 22102 2746
rect 22114 2694 22166 2746
rect 31858 2694 31910 2746
rect 31922 2694 31974 2746
rect 31986 2694 32038 2746
rect 32050 2694 32102 2746
rect 32114 2694 32166 2746
rect 41858 2694 41910 2746
rect 41922 2694 41974 2746
rect 41986 2694 42038 2746
rect 42050 2694 42102 2746
rect 42114 2694 42166 2746
rect 51858 2694 51910 2746
rect 51922 2694 51974 2746
rect 51986 2694 52038 2746
rect 52050 2694 52102 2746
rect 52114 2694 52166 2746
rect 61858 2694 61910 2746
rect 61922 2694 61974 2746
rect 61986 2694 62038 2746
rect 62050 2694 62102 2746
rect 62114 2694 62166 2746
rect 71858 2694 71910 2746
rect 71922 2694 71974 2746
rect 71986 2694 72038 2746
rect 72050 2694 72102 2746
rect 72114 2694 72166 2746
rect 18144 2592 18196 2644
rect 19156 2592 19208 2644
rect 19892 2635 19944 2644
rect 19892 2601 19901 2635
rect 19901 2601 19935 2635
rect 19935 2601 19944 2635
rect 19892 2592 19944 2601
rect 20812 2592 20864 2644
rect 21732 2592 21784 2644
rect 23296 2592 23348 2644
rect 24032 2592 24084 2644
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 25320 2635 25372 2644
rect 25320 2601 25329 2635
rect 25329 2601 25363 2635
rect 25363 2601 25372 2635
rect 25320 2592 25372 2601
rect 27528 2635 27580 2644
rect 27528 2601 27537 2635
rect 27537 2601 27571 2635
rect 27571 2601 27580 2635
rect 27528 2592 27580 2601
rect 29092 2592 29144 2644
rect 31576 2592 31628 2644
rect 33140 2635 33192 2644
rect 33140 2601 33149 2635
rect 33149 2601 33183 2635
rect 33183 2601 33192 2635
rect 33140 2592 33192 2601
rect 34060 2592 34112 2644
rect 36176 2592 36228 2644
rect 46572 2592 46624 2644
rect 48228 2592 48280 2644
rect 53932 2635 53984 2644
rect 53932 2601 53941 2635
rect 53941 2601 53975 2635
rect 53975 2601 53984 2635
rect 53932 2592 53984 2601
rect 60740 2592 60792 2644
rect 67364 2592 67416 2644
rect 16948 2388 17000 2440
rect 25872 2524 25924 2576
rect 30472 2524 30524 2576
rect 19708 2456 19760 2508
rect 20812 2456 20864 2508
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 20260 2388 20312 2440
rect 20628 2320 20680 2372
rect 21364 2388 21416 2440
rect 25964 2456 26016 2508
rect 28448 2456 28500 2508
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 39304 2567 39356 2576
rect 39304 2533 39313 2567
rect 39313 2533 39347 2567
rect 39347 2533 39356 2567
rect 39304 2524 39356 2533
rect 44732 2524 44784 2576
rect 47216 2524 47268 2576
rect 55312 2524 55364 2576
rect 68744 2524 68796 2576
rect 65800 2456 65852 2508
rect 67456 2499 67508 2508
rect 67456 2465 67465 2499
rect 67465 2465 67499 2499
rect 67499 2465 67508 2499
rect 67456 2456 67508 2465
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 24032 2388 24084 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2388 25280 2440
rect 26056 2431 26108 2440
rect 26056 2397 26065 2431
rect 26065 2397 26099 2431
rect 26099 2397 26108 2431
rect 26056 2388 26108 2397
rect 26884 2388 26936 2440
rect 27436 2388 27488 2440
rect 28264 2388 28316 2440
rect 28632 2431 28684 2440
rect 28632 2397 28641 2431
rect 28641 2397 28675 2431
rect 28675 2397 28684 2431
rect 28632 2388 28684 2397
rect 29184 2388 29236 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 32220 2388 32272 2440
rect 32496 2431 32548 2440
rect 32496 2397 32505 2431
rect 32505 2397 32539 2431
rect 32539 2397 32548 2431
rect 32496 2388 32548 2397
rect 33600 2431 33652 2440
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 36544 2431 36596 2440
rect 36544 2397 36553 2431
rect 36553 2397 36587 2431
rect 36587 2397 36596 2431
rect 36544 2388 36596 2397
rect 21732 2320 21784 2372
rect 17776 2252 17828 2304
rect 18328 2252 18380 2304
rect 20904 2252 20956 2304
rect 26700 2295 26752 2304
rect 26700 2261 26709 2295
rect 26709 2261 26743 2295
rect 26743 2261 26752 2295
rect 26700 2252 26752 2261
rect 26792 2295 26844 2304
rect 26792 2261 26801 2295
rect 26801 2261 26835 2295
rect 26835 2261 26844 2295
rect 26792 2252 26844 2261
rect 28540 2295 28592 2304
rect 28540 2261 28549 2295
rect 28549 2261 28583 2295
rect 28583 2261 28592 2295
rect 28540 2252 28592 2261
rect 29092 2252 29144 2304
rect 30288 2295 30340 2304
rect 30288 2261 30297 2295
rect 30297 2261 30331 2295
rect 30331 2261 30340 2295
rect 30288 2252 30340 2261
rect 31300 2252 31352 2304
rect 41420 2388 41472 2440
rect 42340 2388 42392 2440
rect 43444 2388 43496 2440
rect 45560 2431 45612 2440
rect 45560 2397 45569 2431
rect 45569 2397 45603 2431
rect 45603 2397 45612 2431
rect 45560 2388 45612 2397
rect 46204 2431 46256 2440
rect 46204 2397 46213 2431
rect 46213 2397 46247 2431
rect 46247 2397 46256 2431
rect 46204 2388 46256 2397
rect 47308 2388 47360 2440
rect 39120 2320 39172 2372
rect 44640 2320 44692 2372
rect 43536 2252 43588 2304
rect 46848 2252 46900 2304
rect 48872 2388 48924 2440
rect 48964 2388 49016 2440
rect 53840 2388 53892 2440
rect 53932 2388 53984 2440
rect 54024 2320 54076 2372
rect 55036 2320 55088 2372
rect 56692 2320 56744 2372
rect 57336 2431 57388 2440
rect 57336 2397 57345 2431
rect 57345 2397 57379 2431
rect 57379 2397 57388 2431
rect 57336 2388 57388 2397
rect 62304 2431 62356 2440
rect 62304 2397 62313 2431
rect 62313 2397 62347 2431
rect 62347 2397 62356 2431
rect 62304 2388 62356 2397
rect 65524 2388 65576 2440
rect 67272 2388 67324 2440
rect 69940 2431 69992 2440
rect 69940 2397 69949 2431
rect 69949 2397 69983 2431
rect 69983 2397 69992 2431
rect 69940 2388 69992 2397
rect 70492 2388 70544 2440
rect 49424 2252 49476 2304
rect 49516 2252 49568 2304
rect 54760 2295 54812 2304
rect 54760 2261 54769 2295
rect 54769 2261 54803 2295
rect 54803 2261 54812 2295
rect 54760 2252 54812 2261
rect 57888 2252 57940 2304
rect 61016 2363 61068 2372
rect 61016 2329 61025 2363
rect 61025 2329 61059 2363
rect 61059 2329 61068 2363
rect 61016 2320 61068 2329
rect 62948 2295 63000 2304
rect 62948 2261 62957 2295
rect 62957 2261 62991 2295
rect 62991 2261 63000 2295
rect 62948 2252 63000 2261
rect 63592 2320 63644 2372
rect 65156 2252 65208 2304
rect 66076 2252 66128 2304
rect 69388 2252 69440 2304
rect 71044 2252 71096 2304
rect 4210 2150 4262 2202
rect 4274 2150 4326 2202
rect 4338 2150 4390 2202
rect 4402 2150 4454 2202
rect 4466 2150 4518 2202
rect 14210 2150 14262 2202
rect 14274 2150 14326 2202
rect 14338 2150 14390 2202
rect 14402 2150 14454 2202
rect 14466 2150 14518 2202
rect 24210 2150 24262 2202
rect 24274 2150 24326 2202
rect 24338 2150 24390 2202
rect 24402 2150 24454 2202
rect 24466 2150 24518 2202
rect 34210 2150 34262 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 44210 2150 44262 2202
rect 44274 2150 44326 2202
rect 44338 2150 44390 2202
rect 44402 2150 44454 2202
rect 44466 2150 44518 2202
rect 54210 2150 54262 2202
rect 54274 2150 54326 2202
rect 54338 2150 54390 2202
rect 54402 2150 54454 2202
rect 54466 2150 54518 2202
rect 64210 2150 64262 2202
rect 64274 2150 64326 2202
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 74210 2150 74262 2202
rect 74274 2150 74326 2202
rect 74338 2150 74390 2202
rect 74402 2150 74454 2202
rect 74466 2150 74518 2202
rect 17592 2048 17644 2100
rect 18236 2048 18288 2100
rect 18328 1980 18380 2032
rect 21456 2048 21508 2100
rect 24584 2048 24636 2100
rect 19432 1980 19484 2032
rect 26976 2048 27028 2100
rect 16396 1912 16448 1964
rect 18420 1912 18472 1964
rect 22376 1912 22428 1964
rect 24952 1912 25004 1964
rect 25872 1955 25924 1964
rect 25872 1921 25881 1955
rect 25881 1921 25915 1955
rect 25915 1921 25924 1955
rect 25872 1912 25924 1921
rect 26792 1980 26844 2032
rect 28540 1980 28592 2032
rect 32312 2048 32364 2100
rect 32496 2091 32548 2100
rect 32496 2057 32505 2091
rect 32505 2057 32539 2091
rect 32539 2057 32548 2091
rect 32496 2048 32548 2057
rect 34612 2091 34664 2100
rect 34612 2057 34621 2091
rect 34621 2057 34655 2091
rect 34655 2057 34664 2091
rect 34612 2048 34664 2057
rect 34704 2048 34756 2100
rect 36176 2048 36228 2100
rect 36728 2048 36780 2100
rect 39120 2091 39172 2100
rect 39120 2057 39129 2091
rect 39129 2057 39163 2091
rect 39163 2057 39172 2091
rect 39120 2048 39172 2057
rect 39304 2048 39356 2100
rect 41696 2048 41748 2100
rect 42248 2048 42300 2100
rect 44824 2048 44876 2100
rect 45468 2048 45520 2100
rect 50436 2048 50488 2100
rect 51540 2048 51592 2100
rect 55036 2091 55088 2100
rect 55036 2057 55045 2091
rect 55045 2057 55079 2091
rect 55079 2057 55088 2091
rect 55036 2048 55088 2057
rect 61108 2048 61160 2100
rect 63592 2091 63644 2100
rect 63592 2057 63601 2091
rect 63601 2057 63635 2091
rect 63635 2057 63644 2091
rect 63592 2048 63644 2057
rect 26700 1912 26752 1964
rect 18052 1844 18104 1896
rect 19340 1844 19392 1896
rect 23204 1887 23256 1896
rect 23204 1853 23213 1887
rect 23213 1853 23247 1887
rect 23247 1853 23256 1887
rect 23204 1844 23256 1853
rect 24676 1844 24728 1896
rect 28448 1844 28500 1896
rect 28816 1844 28868 1896
rect 29092 1955 29144 1964
rect 29092 1921 29101 1955
rect 29101 1921 29135 1955
rect 29135 1921 29144 1955
rect 29092 1912 29144 1921
rect 29552 1912 29604 1964
rect 66904 1980 66956 2032
rect 67272 2091 67324 2100
rect 67272 2057 67281 2091
rect 67281 2057 67315 2091
rect 67315 2057 67324 2091
rect 67272 2048 67324 2057
rect 67916 1980 67968 2032
rect 69204 1980 69256 2032
rect 70124 1980 70176 2032
rect 29920 1912 29972 1964
rect 30288 1844 30340 1896
rect 31300 1955 31352 1964
rect 31300 1921 31309 1955
rect 31309 1921 31343 1955
rect 31343 1921 31352 1955
rect 31300 1912 31352 1921
rect 34060 1912 34112 1964
rect 34796 1955 34848 1964
rect 34796 1921 34805 1955
rect 34805 1921 34839 1955
rect 34839 1921 34848 1955
rect 34796 1912 34848 1921
rect 39028 1912 39080 1964
rect 42892 1912 42944 1964
rect 42984 1955 43036 1964
rect 42984 1921 42993 1955
rect 42993 1921 43027 1955
rect 43027 1921 43036 1955
rect 42984 1912 43036 1921
rect 32404 1844 32456 1896
rect 34612 1844 34664 1896
rect 36176 1887 36228 1896
rect 36176 1853 36185 1887
rect 36185 1853 36219 1887
rect 36219 1853 36228 1887
rect 36176 1844 36228 1853
rect 37556 1887 37608 1896
rect 37556 1853 37565 1887
rect 37565 1853 37599 1887
rect 37599 1853 37608 1887
rect 37556 1844 37608 1853
rect 41144 1887 41196 1896
rect 41144 1853 41153 1887
rect 41153 1853 41187 1887
rect 41187 1853 41196 1887
rect 41144 1844 41196 1853
rect 35900 1776 35952 1828
rect 35992 1776 36044 1828
rect 41512 1776 41564 1828
rect 42984 1776 43036 1828
rect 45652 1912 45704 1964
rect 46848 1912 46900 1964
rect 47584 1912 47636 1964
rect 49516 1955 49568 1964
rect 49516 1921 49525 1955
rect 49525 1921 49559 1955
rect 49559 1921 49568 1955
rect 49516 1912 49568 1921
rect 53104 1955 53156 1964
rect 53104 1921 53113 1955
rect 53113 1921 53147 1955
rect 53147 1921 53156 1955
rect 53104 1912 53156 1921
rect 54760 1912 54812 1964
rect 56416 1955 56468 1964
rect 56416 1921 56425 1955
rect 56425 1921 56459 1955
rect 56459 1921 56468 1955
rect 56416 1912 56468 1921
rect 57888 1955 57940 1964
rect 57888 1921 57897 1955
rect 57897 1921 57931 1955
rect 57931 1921 57940 1955
rect 57888 1912 57940 1921
rect 61384 1955 61436 1964
rect 61384 1921 61393 1955
rect 61393 1921 61427 1955
rect 61427 1921 61436 1955
rect 61384 1912 61436 1921
rect 62948 1955 63000 1964
rect 62948 1921 62957 1955
rect 62957 1921 62991 1955
rect 62991 1921 63000 1955
rect 62948 1912 63000 1921
rect 64604 1955 64656 1964
rect 64604 1921 64613 1955
rect 64613 1921 64647 1955
rect 64647 1921 64656 1955
rect 64604 1912 64656 1921
rect 66076 1955 66128 1964
rect 66076 1921 66085 1955
rect 66085 1921 66119 1955
rect 66119 1921 66128 1955
rect 66076 1912 66128 1921
rect 67180 1912 67232 1964
rect 69388 1955 69440 1964
rect 69388 1921 69397 1955
rect 69397 1921 69431 1955
rect 69431 1921 69440 1955
rect 69388 1912 69440 1921
rect 69664 1955 69716 1964
rect 69664 1921 69673 1955
rect 69673 1921 69707 1955
rect 69707 1921 69716 1955
rect 69664 1912 69716 1921
rect 71044 1955 71096 1964
rect 71044 1921 71053 1955
rect 71053 1921 71087 1955
rect 71087 1921 71096 1955
rect 71044 1912 71096 1921
rect 46020 1887 46072 1896
rect 46020 1853 46029 1887
rect 46029 1853 46063 1887
rect 46063 1853 46072 1887
rect 46020 1844 46072 1853
rect 46204 1887 46256 1896
rect 46204 1853 46213 1887
rect 46213 1853 46247 1887
rect 46247 1853 46256 1887
rect 46204 1844 46256 1853
rect 47860 1844 47912 1896
rect 51264 1887 51316 1896
rect 51264 1853 51273 1887
rect 51273 1853 51307 1887
rect 51307 1853 51316 1887
rect 51264 1844 51316 1853
rect 52828 1844 52880 1896
rect 55588 1887 55640 1896
rect 55588 1853 55597 1887
rect 55597 1853 55631 1887
rect 55631 1853 55640 1887
rect 55588 1844 55640 1853
rect 56140 1844 56192 1896
rect 59360 1844 59412 1896
rect 60556 1887 60608 1896
rect 60556 1853 60565 1887
rect 60565 1853 60599 1887
rect 60599 1853 60608 1887
rect 60556 1844 60608 1853
rect 61108 1844 61160 1896
rect 63868 1887 63920 1896
rect 63868 1853 63877 1887
rect 63877 1853 63911 1887
rect 63911 1853 63920 1887
rect 63868 1844 63920 1853
rect 64696 1844 64748 1896
rect 72240 1844 72292 1896
rect 46940 1776 46992 1828
rect 23388 1708 23440 1760
rect 29000 1708 29052 1760
rect 34704 1708 34756 1760
rect 38568 1751 38620 1760
rect 38568 1717 38577 1751
rect 38577 1717 38611 1751
rect 38611 1717 38620 1751
rect 38568 1708 38620 1717
rect 47216 1708 47268 1760
rect 55772 1776 55824 1828
rect 65432 1776 65484 1828
rect 69388 1776 69440 1828
rect 53380 1708 53432 1760
rect 57244 1708 57296 1760
rect 62396 1708 62448 1760
rect 65156 1708 65208 1760
rect 73160 1708 73212 1760
rect 1858 1606 1910 1658
rect 1922 1606 1974 1658
rect 1986 1606 2038 1658
rect 2050 1606 2102 1658
rect 2114 1606 2166 1658
rect 11858 1606 11910 1658
rect 11922 1606 11974 1658
rect 11986 1606 12038 1658
rect 12050 1606 12102 1658
rect 12114 1606 12166 1658
rect 21858 1606 21910 1658
rect 21922 1606 21974 1658
rect 21986 1606 22038 1658
rect 22050 1606 22102 1658
rect 22114 1606 22166 1658
rect 31858 1606 31910 1658
rect 31922 1606 31974 1658
rect 31986 1606 32038 1658
rect 32050 1606 32102 1658
rect 32114 1606 32166 1658
rect 41858 1606 41910 1658
rect 41922 1606 41974 1658
rect 41986 1606 42038 1658
rect 42050 1606 42102 1658
rect 42114 1606 42166 1658
rect 51858 1606 51910 1658
rect 51922 1606 51974 1658
rect 51986 1606 52038 1658
rect 52050 1606 52102 1658
rect 52114 1606 52166 1658
rect 61858 1606 61910 1658
rect 61922 1606 61974 1658
rect 61986 1606 62038 1658
rect 62050 1606 62102 1658
rect 62114 1606 62166 1658
rect 71858 1606 71910 1658
rect 71922 1606 71974 1658
rect 71986 1606 72038 1658
rect 72050 1606 72102 1658
rect 72114 1606 72166 1658
rect 22928 1504 22980 1556
rect 26056 1504 26108 1556
rect 28632 1504 28684 1556
rect 31024 1504 31076 1556
rect 37556 1504 37608 1556
rect 41144 1504 41196 1556
rect 31116 1436 31168 1488
rect 35164 1436 35216 1488
rect 36544 1436 36596 1488
rect 38568 1436 38620 1488
rect 45468 1504 45520 1556
rect 45560 1504 45612 1556
rect 46940 1504 46992 1556
rect 51264 1504 51316 1556
rect 61016 1504 61068 1556
rect 63868 1504 63920 1556
rect 69940 1504 69992 1556
rect 41696 1436 41748 1488
rect 47032 1436 47084 1488
rect 27988 1368 28040 1420
rect 28448 1368 28500 1420
rect 35072 1368 35124 1420
rect 37924 1368 37976 1420
rect 41236 1368 41288 1420
rect 5080 1343 5132 1352
rect 5080 1309 5089 1343
rect 5089 1309 5123 1343
rect 5123 1309 5132 1343
rect 5080 1300 5132 1309
rect 15292 1300 15344 1352
rect 17500 1300 17552 1352
rect 17776 1343 17828 1352
rect 17776 1309 17785 1343
rect 17785 1309 17819 1343
rect 17819 1309 17828 1343
rect 17776 1300 17828 1309
rect 3148 1232 3200 1284
rect 15936 1232 15988 1284
rect 15568 1207 15620 1216
rect 15568 1173 15577 1207
rect 15577 1173 15611 1207
rect 15611 1173 15620 1207
rect 15568 1164 15620 1173
rect 19064 1300 19116 1352
rect 19432 1275 19484 1284
rect 19432 1241 19441 1275
rect 19441 1241 19475 1275
rect 19475 1241 19484 1275
rect 19432 1232 19484 1241
rect 19800 1343 19852 1352
rect 19800 1309 19809 1343
rect 19809 1309 19843 1343
rect 19843 1309 19852 1343
rect 19800 1300 19852 1309
rect 22560 1300 22612 1352
rect 22284 1232 22336 1284
rect 23572 1232 23624 1284
rect 26332 1300 26384 1352
rect 25780 1275 25832 1284
rect 25780 1241 25789 1275
rect 25789 1241 25823 1275
rect 25823 1241 25832 1275
rect 25780 1232 25832 1241
rect 26516 1164 26568 1216
rect 28080 1343 28132 1352
rect 28080 1309 28089 1343
rect 28089 1309 28123 1343
rect 28123 1309 28132 1343
rect 28080 1300 28132 1309
rect 29460 1343 29512 1352
rect 29460 1309 29469 1343
rect 29469 1309 29503 1343
rect 29503 1309 29512 1343
rect 29460 1300 29512 1309
rect 30380 1300 30432 1352
rect 28540 1232 28592 1284
rect 32864 1300 32916 1352
rect 33232 1343 33284 1352
rect 33232 1309 33241 1343
rect 33241 1309 33275 1343
rect 33275 1309 33284 1343
rect 33232 1300 33284 1309
rect 27896 1164 27948 1216
rect 31300 1232 31352 1284
rect 33048 1232 33100 1284
rect 33600 1164 33652 1216
rect 35624 1343 35676 1352
rect 35624 1309 35633 1343
rect 35633 1309 35667 1343
rect 35667 1309 35676 1343
rect 35624 1300 35676 1309
rect 37372 1343 37424 1352
rect 37372 1309 37381 1343
rect 37381 1309 37415 1343
rect 37415 1309 37424 1343
rect 37372 1300 37424 1309
rect 38016 1343 38068 1352
rect 38016 1309 38025 1343
rect 38025 1309 38059 1343
rect 38059 1309 38068 1343
rect 38016 1300 38068 1309
rect 39764 1343 39816 1352
rect 39764 1309 39773 1343
rect 39773 1309 39807 1343
rect 39807 1309 39816 1343
rect 39764 1300 39816 1309
rect 40776 1300 40828 1352
rect 42432 1343 42484 1352
rect 42432 1309 42441 1343
rect 42441 1309 42475 1343
rect 42475 1309 42484 1343
rect 42432 1300 42484 1309
rect 42892 1300 42944 1352
rect 44640 1368 44692 1420
rect 44824 1368 44876 1420
rect 46204 1368 46256 1420
rect 49608 1368 49660 1420
rect 59452 1368 59504 1420
rect 62764 1368 62816 1420
rect 67732 1368 67784 1420
rect 71044 1368 71096 1420
rect 44732 1300 44784 1352
rect 44916 1343 44968 1352
rect 44916 1309 44925 1343
rect 44925 1309 44959 1343
rect 44959 1309 44968 1343
rect 44916 1300 44968 1309
rect 36176 1232 36228 1284
rect 36268 1232 36320 1284
rect 39580 1232 39632 1284
rect 43996 1232 44048 1284
rect 45100 1232 45152 1284
rect 47492 1343 47544 1352
rect 47492 1309 47501 1343
rect 47501 1309 47535 1343
rect 47535 1309 47544 1343
rect 47492 1300 47544 1309
rect 48872 1300 48924 1352
rect 49424 1300 49476 1352
rect 50068 1343 50120 1352
rect 50068 1309 50077 1343
rect 50077 1309 50111 1343
rect 50111 1309 50120 1343
rect 50068 1300 50120 1309
rect 50620 1300 50672 1352
rect 52644 1343 52696 1352
rect 52644 1309 52653 1343
rect 52653 1309 52687 1343
rect 52687 1309 52696 1343
rect 52644 1300 52696 1309
rect 53840 1300 53892 1352
rect 51172 1232 51224 1284
rect 35716 1164 35768 1216
rect 46020 1164 46072 1216
rect 52276 1164 52328 1216
rect 55220 1343 55272 1352
rect 55220 1309 55229 1343
rect 55229 1309 55263 1343
rect 55263 1309 55272 1343
rect 55220 1300 55272 1309
rect 56692 1343 56744 1352
rect 56692 1309 56701 1343
rect 56701 1309 56735 1343
rect 56735 1309 56744 1343
rect 56692 1300 56744 1309
rect 57244 1343 57296 1352
rect 57244 1309 57253 1343
rect 57253 1309 57287 1343
rect 57287 1309 57296 1343
rect 57244 1300 57296 1309
rect 57980 1343 58032 1352
rect 57980 1309 57989 1343
rect 57989 1309 58023 1343
rect 58023 1309 58032 1343
rect 57980 1300 58032 1309
rect 59360 1343 59412 1352
rect 59360 1309 59369 1343
rect 59369 1309 59403 1343
rect 59403 1309 59412 1343
rect 59360 1300 59412 1309
rect 54576 1232 54628 1284
rect 57796 1232 57848 1284
rect 58900 1232 58952 1284
rect 60372 1343 60424 1352
rect 60372 1309 60381 1343
rect 60381 1309 60415 1343
rect 60415 1309 60424 1343
rect 60372 1300 60424 1309
rect 62396 1343 62448 1352
rect 62396 1309 62405 1343
rect 62405 1309 62439 1343
rect 62439 1309 62448 1343
rect 62396 1300 62448 1309
rect 63040 1343 63092 1352
rect 63040 1309 63049 1343
rect 63049 1309 63083 1343
rect 63083 1309 63092 1343
rect 63040 1300 63092 1309
rect 63868 1300 63920 1352
rect 65156 1300 65208 1352
rect 66260 1343 66312 1352
rect 66260 1309 66269 1343
rect 66269 1309 66303 1343
rect 66303 1309 66312 1343
rect 66260 1300 66312 1309
rect 68284 1343 68336 1352
rect 68284 1309 68293 1343
rect 68293 1309 68327 1343
rect 68327 1309 68336 1343
rect 68284 1300 68336 1309
rect 68836 1300 68888 1352
rect 71228 1343 71280 1352
rect 71228 1309 71237 1343
rect 71237 1309 71271 1343
rect 71271 1309 71280 1343
rect 71228 1300 71280 1309
rect 73160 1300 73212 1352
rect 73252 1343 73304 1352
rect 73252 1309 73261 1343
rect 73261 1309 73295 1343
rect 73295 1309 73304 1343
rect 73252 1300 73304 1309
rect 66076 1232 66128 1284
rect 70032 1232 70084 1284
rect 67364 1164 67416 1216
rect 72700 1164 72752 1216
rect 4210 1062 4262 1114
rect 4274 1062 4326 1114
rect 4338 1062 4390 1114
rect 4402 1062 4454 1114
rect 4466 1062 4518 1114
rect 14210 1062 14262 1114
rect 14274 1062 14326 1114
rect 14338 1062 14390 1114
rect 14402 1062 14454 1114
rect 14466 1062 14518 1114
rect 24210 1062 24262 1114
rect 24274 1062 24326 1114
rect 24338 1062 24390 1114
rect 24402 1062 24454 1114
rect 24466 1062 24518 1114
rect 34210 1062 34262 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 44210 1062 44262 1114
rect 44274 1062 44326 1114
rect 44338 1062 44390 1114
rect 44402 1062 44454 1114
rect 44466 1062 44518 1114
rect 54210 1062 54262 1114
rect 54274 1062 54326 1114
rect 54338 1062 54390 1114
rect 54402 1062 54454 1114
rect 54466 1062 54518 1114
rect 64210 1062 64262 1114
rect 64274 1062 64326 1114
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 74210 1062 74262 1114
rect 74274 1062 74326 1114
rect 74338 1062 74390 1114
rect 74402 1062 74454 1114
rect 74466 1062 74518 1114
rect 5080 960 5132 1012
rect 23940 960 23992 1012
rect 31392 960 31444 1012
rect 35624 960 35676 1012
rect 15568 892 15620 944
rect 20720 892 20772 944
rect 32864 892 32916 944
rect 33508 892 33560 944
rect 19432 824 19484 876
rect 43812 824 43864 876
<< metal2 >>
rect 71836 85434 72188 86000
rect 71836 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 72188 85434
rect 2020 84588 2124 84616
rect 2020 84532 2044 84588
rect 2100 84532 2124 84588
rect 2020 84508 2124 84532
rect 2020 84452 2044 84508
rect 2100 84452 2124 84508
rect 2020 84428 2124 84452
rect 2020 84372 2044 84428
rect 2100 84372 2124 84428
rect 2020 84348 2124 84372
rect 2020 84292 2044 84348
rect 2100 84292 2124 84348
rect 2020 84264 2124 84292
rect 5521 84588 5615 84616
rect 5521 84532 5540 84588
rect 5596 84532 5615 84588
rect 5521 84508 5615 84532
rect 5521 84452 5540 84508
rect 5596 84452 5615 84508
rect 5521 84428 5615 84452
rect 5521 84372 5540 84428
rect 5596 84372 5615 84428
rect 5521 84348 5615 84372
rect 5521 84292 5540 84348
rect 5596 84292 5615 84348
rect 5521 84264 5615 84292
rect 8411 84588 8505 84616
rect 8411 84532 8430 84588
rect 8486 84532 8505 84588
rect 8411 84508 8505 84532
rect 8411 84452 8430 84508
rect 8486 84452 8505 84508
rect 8411 84428 8505 84452
rect 8411 84372 8430 84428
rect 8486 84372 8505 84428
rect 8411 84348 8505 84372
rect 8411 84292 8430 84348
rect 8486 84292 8505 84348
rect 8411 84264 8505 84292
rect 11301 84588 11395 84616
rect 11301 84532 11320 84588
rect 11376 84532 11395 84588
rect 11301 84508 11395 84532
rect 11301 84452 11320 84508
rect 11376 84452 11395 84508
rect 11301 84428 11395 84452
rect 11301 84372 11320 84428
rect 11376 84372 11395 84428
rect 11301 84348 11395 84372
rect 11301 84292 11320 84348
rect 11376 84292 11395 84348
rect 11301 84264 11395 84292
rect 14191 84588 14285 84616
rect 14191 84532 14210 84588
rect 14266 84532 14285 84588
rect 14191 84508 14285 84532
rect 14191 84452 14210 84508
rect 14266 84452 14285 84508
rect 14191 84428 14285 84452
rect 14191 84372 14210 84428
rect 14266 84372 14285 84428
rect 14191 84348 14285 84372
rect 14191 84292 14210 84348
rect 14266 84292 14285 84348
rect 14191 84264 14285 84292
rect 17081 84588 17175 84616
rect 17081 84532 17100 84588
rect 17156 84532 17175 84588
rect 17081 84508 17175 84532
rect 17081 84452 17100 84508
rect 17156 84452 17175 84508
rect 17081 84428 17175 84452
rect 17081 84372 17100 84428
rect 17156 84372 17175 84428
rect 17081 84348 17175 84372
rect 17081 84292 17100 84348
rect 17156 84292 17175 84348
rect 17081 84264 17175 84292
rect 19971 84588 20065 84616
rect 19971 84532 19990 84588
rect 20046 84532 20065 84588
rect 19971 84508 20065 84532
rect 19971 84452 19990 84508
rect 20046 84452 20065 84508
rect 19971 84428 20065 84452
rect 19971 84372 19990 84428
rect 20046 84372 20065 84428
rect 19971 84348 20065 84372
rect 19971 84292 19990 84348
rect 20046 84292 20065 84348
rect 19971 84264 20065 84292
rect 22861 84588 22955 84616
rect 22861 84532 22880 84588
rect 22936 84532 22955 84588
rect 22861 84508 22955 84532
rect 22861 84452 22880 84508
rect 22936 84452 22955 84508
rect 22861 84428 22955 84452
rect 22861 84372 22880 84428
rect 22936 84372 22955 84428
rect 22861 84348 22955 84372
rect 22861 84292 22880 84348
rect 22936 84292 22955 84348
rect 22861 84264 22955 84292
rect 25751 84588 25845 84616
rect 25751 84532 25770 84588
rect 25826 84532 25845 84588
rect 25751 84508 25845 84532
rect 25751 84452 25770 84508
rect 25826 84452 25845 84508
rect 25751 84428 25845 84452
rect 25751 84372 25770 84428
rect 25826 84372 25845 84428
rect 25751 84348 25845 84372
rect 25751 84292 25770 84348
rect 25826 84292 25845 84348
rect 25751 84264 25845 84292
rect 28641 84588 28735 84616
rect 28641 84532 28660 84588
rect 28716 84532 28735 84588
rect 28641 84508 28735 84532
rect 28641 84452 28660 84508
rect 28716 84452 28735 84508
rect 28641 84428 28735 84452
rect 28641 84372 28660 84428
rect 28716 84372 28735 84428
rect 28641 84348 28735 84372
rect 28641 84292 28660 84348
rect 28716 84292 28735 84348
rect 28641 84264 28735 84292
rect 31531 84588 31625 84616
rect 31531 84532 31550 84588
rect 31606 84532 31625 84588
rect 31531 84508 31625 84532
rect 31531 84452 31550 84508
rect 31606 84452 31625 84508
rect 31531 84428 31625 84452
rect 31531 84372 31550 84428
rect 31606 84372 31625 84428
rect 31531 84348 31625 84372
rect 31531 84292 31550 84348
rect 31606 84292 31625 84348
rect 31531 84264 31625 84292
rect 34421 84588 34515 84616
rect 34421 84532 34440 84588
rect 34496 84532 34515 84588
rect 34421 84508 34515 84532
rect 34421 84452 34440 84508
rect 34496 84452 34515 84508
rect 34421 84428 34515 84452
rect 34421 84372 34440 84428
rect 34496 84372 34515 84428
rect 34421 84348 34515 84372
rect 34421 84292 34440 84348
rect 34496 84292 34515 84348
rect 34421 84264 34515 84292
rect 37311 84588 37405 84616
rect 37311 84532 37330 84588
rect 37386 84532 37405 84588
rect 37311 84508 37405 84532
rect 37311 84452 37330 84508
rect 37386 84452 37405 84508
rect 37311 84428 37405 84452
rect 37311 84372 37330 84428
rect 37386 84372 37405 84428
rect 37311 84348 37405 84372
rect 37311 84292 37330 84348
rect 37386 84292 37405 84348
rect 37311 84264 37405 84292
rect 40201 84588 40295 84616
rect 40201 84532 40220 84588
rect 40276 84532 40295 84588
rect 40201 84508 40295 84532
rect 40201 84452 40220 84508
rect 40276 84452 40295 84508
rect 40201 84428 40295 84452
rect 40201 84372 40220 84428
rect 40276 84372 40295 84428
rect 40201 84348 40295 84372
rect 40201 84292 40220 84348
rect 40276 84292 40295 84348
rect 40201 84264 40295 84292
rect 43091 84588 43185 84616
rect 43091 84532 43110 84588
rect 43166 84532 43185 84588
rect 43091 84508 43185 84532
rect 43091 84452 43110 84508
rect 43166 84452 43185 84508
rect 43091 84428 43185 84452
rect 43091 84372 43110 84428
rect 43166 84372 43185 84428
rect 43091 84348 43185 84372
rect 43091 84292 43110 84348
rect 43166 84292 43185 84348
rect 43091 84264 43185 84292
rect 45981 84588 46075 84616
rect 45981 84532 46000 84588
rect 46056 84532 46075 84588
rect 45981 84508 46075 84532
rect 45981 84452 46000 84508
rect 46056 84452 46075 84508
rect 45981 84428 46075 84452
rect 45981 84372 46000 84428
rect 46056 84372 46075 84428
rect 45981 84348 46075 84372
rect 45981 84292 46000 84348
rect 46056 84292 46075 84348
rect 45981 84264 46075 84292
rect 48989 84588 49083 84616
rect 48989 84532 49008 84588
rect 49064 84532 49083 84588
rect 48989 84508 49083 84532
rect 48989 84452 49008 84508
rect 49064 84452 49083 84508
rect 48989 84428 49083 84452
rect 48989 84372 49008 84428
rect 49064 84372 49083 84428
rect 48989 84348 49083 84372
rect 48989 84292 49008 84348
rect 49064 84292 49083 84348
rect 48989 84264 49083 84292
rect 52210 84588 52320 84616
rect 52210 84532 52237 84588
rect 52293 84532 52320 84588
rect 52210 84508 52320 84532
rect 52210 84452 52237 84508
rect 52293 84452 52320 84508
rect 52210 84428 52320 84452
rect 52210 84372 52237 84428
rect 52293 84372 52320 84428
rect 52210 84348 52320 84372
rect 52210 84292 52237 84348
rect 52293 84292 52320 84348
rect 52210 84264 52320 84292
rect 53602 84588 53730 84616
rect 53602 84532 53638 84588
rect 53694 84532 53730 84588
rect 53602 84508 53730 84532
rect 53602 84452 53638 84508
rect 53694 84452 53730 84508
rect 53602 84428 53730 84452
rect 53602 84372 53638 84428
rect 53694 84372 53730 84428
rect 53602 84348 53730 84372
rect 53602 84292 53638 84348
rect 53694 84292 53730 84348
rect 53602 84264 53730 84292
rect 53770 84588 53898 84616
rect 53770 84532 53806 84588
rect 53862 84532 53898 84588
rect 53770 84508 53898 84532
rect 53770 84452 53806 84508
rect 53862 84452 53898 84508
rect 53770 84428 53898 84452
rect 53770 84372 53806 84428
rect 53862 84372 53898 84428
rect 53770 84348 53898 84372
rect 53770 84292 53806 84348
rect 53862 84292 53898 84348
rect 53770 84264 53898 84292
rect 54514 84588 54642 84616
rect 54514 84532 54550 84588
rect 54606 84532 54642 84588
rect 54514 84508 54642 84532
rect 54514 84452 54550 84508
rect 54606 84452 54642 84508
rect 54514 84428 54642 84452
rect 54514 84372 54550 84428
rect 54606 84372 54642 84428
rect 54514 84348 54642 84372
rect 54514 84292 54550 84348
rect 54606 84292 54642 84348
rect 54514 84264 54642 84292
rect 54910 84588 55026 84616
rect 54910 84532 54940 84588
rect 54996 84532 55026 84588
rect 54910 84508 55026 84532
rect 54910 84452 54940 84508
rect 54996 84452 55026 84508
rect 54910 84428 55026 84452
rect 54910 84372 54940 84428
rect 54996 84372 55026 84428
rect 54910 84348 55026 84372
rect 54910 84292 54940 84348
rect 54996 84292 55026 84348
rect 54910 84264 55026 84292
rect 55620 84588 55748 84616
rect 55620 84532 55656 84588
rect 55712 84532 55748 84588
rect 55620 84508 55748 84532
rect 55620 84452 55656 84508
rect 55712 84452 55748 84508
rect 55620 84428 55748 84452
rect 55620 84372 55656 84428
rect 55712 84372 55748 84428
rect 55620 84348 55748 84372
rect 55620 84292 55656 84348
rect 55712 84292 55748 84348
rect 55620 84264 55748 84292
rect 56198 84588 56326 84616
rect 56198 84532 56234 84588
rect 56290 84532 56326 84588
rect 56198 84508 56326 84532
rect 56198 84452 56234 84508
rect 56290 84452 56326 84508
rect 56198 84428 56326 84452
rect 56198 84372 56234 84428
rect 56290 84372 56326 84428
rect 56198 84348 56326 84372
rect 56198 84292 56234 84348
rect 56290 84292 56326 84348
rect 56198 84264 56326 84292
rect 56649 84588 56765 84616
rect 56649 84532 56679 84588
rect 56735 84532 56765 84588
rect 56649 84508 56765 84532
rect 56649 84452 56679 84508
rect 56735 84452 56765 84508
rect 56649 84428 56765 84452
rect 56649 84372 56679 84428
rect 56735 84372 56765 84428
rect 56649 84348 56765 84372
rect 56649 84292 56679 84348
rect 56735 84292 56765 84348
rect 56649 84264 56765 84292
rect 56953 84588 57069 84616
rect 56953 84532 56983 84588
rect 57039 84532 57069 84588
rect 56953 84508 57069 84532
rect 56953 84452 56983 84508
rect 57039 84452 57069 84508
rect 56953 84428 57069 84452
rect 56953 84372 56983 84428
rect 57039 84372 57069 84428
rect 56953 84348 57069 84372
rect 56953 84292 56983 84348
rect 57039 84292 57069 84348
rect 56953 84264 57069 84292
rect 57795 84588 57911 84616
rect 57795 84532 57825 84588
rect 57881 84532 57911 84588
rect 57795 84508 57911 84532
rect 57795 84452 57825 84508
rect 57881 84452 57911 84508
rect 57795 84428 57911 84452
rect 57795 84372 57825 84428
rect 57881 84372 57911 84428
rect 57795 84348 57911 84372
rect 57795 84292 57825 84348
rect 57881 84292 57911 84348
rect 57795 84264 57911 84292
rect 58461 84588 58525 84616
rect 58461 84532 58465 84588
rect 58521 84532 58525 84588
rect 58461 84508 58525 84532
rect 58461 84452 58465 84508
rect 58521 84452 58525 84508
rect 58461 84428 58525 84452
rect 58461 84372 58465 84428
rect 58521 84372 58525 84428
rect 58461 84348 58525 84372
rect 58461 84292 58465 84348
rect 58521 84292 58525 84348
rect 58461 84264 58525 84292
rect 59018 84588 59134 84616
rect 59018 84532 59048 84588
rect 59104 84532 59134 84588
rect 59018 84508 59134 84532
rect 59018 84452 59048 84508
rect 59104 84452 59134 84508
rect 59018 84428 59134 84452
rect 59018 84372 59048 84428
rect 59104 84372 59134 84428
rect 59018 84348 59134 84372
rect 59018 84292 59048 84348
rect 59104 84292 59134 84348
rect 59018 84264 59134 84292
rect 60296 84588 60412 84616
rect 60296 84532 60326 84588
rect 60382 84532 60412 84588
rect 60296 84508 60412 84532
rect 60296 84452 60326 84508
rect 60382 84452 60412 84508
rect 60296 84428 60412 84452
rect 60296 84372 60326 84428
rect 60382 84372 60412 84428
rect 60296 84348 60412 84372
rect 60296 84292 60326 84348
rect 60382 84292 60412 84348
rect 60296 84264 60412 84292
rect 60454 84588 60570 84616
rect 60454 84532 60484 84588
rect 60540 84532 60570 84588
rect 60454 84508 60570 84532
rect 60454 84452 60484 84508
rect 60540 84452 60570 84508
rect 60454 84428 60570 84452
rect 60454 84372 60484 84428
rect 60540 84372 60570 84428
rect 60454 84348 60570 84372
rect 60454 84292 60484 84348
rect 60540 84292 60570 84348
rect 60454 84264 60570 84292
rect 62509 84588 62683 84616
rect 62509 84532 62528 84588
rect 62584 84532 62608 84588
rect 62664 84532 62683 84588
rect 62509 84508 62683 84532
rect 62509 84452 62528 84508
rect 62584 84452 62608 84508
rect 62664 84452 62683 84508
rect 62509 84428 62683 84452
rect 62509 84372 62528 84428
rect 62584 84372 62608 84428
rect 62664 84372 62683 84428
rect 62509 84348 62683 84372
rect 62509 84292 62528 84348
rect 62584 84292 62608 84348
rect 62664 84292 62683 84348
rect 62509 84264 62683 84292
rect 71836 84346 72188 85382
rect 71836 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 72188 84346
rect 64880 84244 64932 84250
rect 64880 84186 64932 84192
rect 2152 82236 2352 82264
rect 2152 82180 2184 82236
rect 2240 82180 2264 82236
rect 2320 82180 2352 82236
rect 2152 82156 2352 82180
rect 2152 82100 2184 82156
rect 2240 82100 2264 82156
rect 2320 82100 2352 82156
rect 2152 82076 2352 82100
rect 2152 82020 2184 82076
rect 2240 82020 2264 82076
rect 2320 82020 2352 82076
rect 2152 81996 2352 82020
rect 2152 81940 2184 81996
rect 2240 81940 2264 81996
rect 2320 81940 2352 81996
rect 2152 81912 2352 81940
rect 5374 82236 5468 82264
rect 5374 82180 5393 82236
rect 5449 82180 5468 82236
rect 5374 82156 5468 82180
rect 5374 82100 5393 82156
rect 5449 82100 5468 82156
rect 5374 82076 5468 82100
rect 5374 82020 5393 82076
rect 5449 82020 5468 82076
rect 5374 81996 5468 82020
rect 5374 81940 5393 81996
rect 5449 81940 5468 81996
rect 5374 81912 5468 81940
rect 8264 82236 8358 82264
rect 8264 82180 8283 82236
rect 8339 82180 8358 82236
rect 8264 82156 8358 82180
rect 8264 82100 8283 82156
rect 8339 82100 8358 82156
rect 8264 82076 8358 82100
rect 8264 82020 8283 82076
rect 8339 82020 8358 82076
rect 8264 81996 8358 82020
rect 8264 81940 8283 81996
rect 8339 81940 8358 81996
rect 8264 81912 8358 81940
rect 11154 82236 11248 82264
rect 11154 82180 11173 82236
rect 11229 82180 11248 82236
rect 11154 82156 11248 82180
rect 11154 82100 11173 82156
rect 11229 82100 11248 82156
rect 11154 82076 11248 82100
rect 11154 82020 11173 82076
rect 11229 82020 11248 82076
rect 11154 81996 11248 82020
rect 11154 81940 11173 81996
rect 11229 81940 11248 81996
rect 11154 81912 11248 81940
rect 14044 82236 14138 82264
rect 14044 82180 14063 82236
rect 14119 82180 14138 82236
rect 14044 82156 14138 82180
rect 14044 82100 14063 82156
rect 14119 82100 14138 82156
rect 14044 82076 14138 82100
rect 14044 82020 14063 82076
rect 14119 82020 14138 82076
rect 14044 81996 14138 82020
rect 14044 81940 14063 81996
rect 14119 81940 14138 81996
rect 14044 81912 14138 81940
rect 16934 82236 17028 82264
rect 16934 82180 16953 82236
rect 17009 82180 17028 82236
rect 16934 82156 17028 82180
rect 16934 82100 16953 82156
rect 17009 82100 17028 82156
rect 16934 82076 17028 82100
rect 16934 82020 16953 82076
rect 17009 82020 17028 82076
rect 16934 81996 17028 82020
rect 16934 81940 16953 81996
rect 17009 81940 17028 81996
rect 16934 81912 17028 81940
rect 19824 82236 19918 82264
rect 19824 82180 19843 82236
rect 19899 82180 19918 82236
rect 19824 82156 19918 82180
rect 19824 82100 19843 82156
rect 19899 82100 19918 82156
rect 19824 82076 19918 82100
rect 19824 82020 19843 82076
rect 19899 82020 19918 82076
rect 19824 81996 19918 82020
rect 19824 81940 19843 81996
rect 19899 81940 19918 81996
rect 19824 81912 19918 81940
rect 22714 82236 22808 82264
rect 22714 82180 22733 82236
rect 22789 82180 22808 82236
rect 22714 82156 22808 82180
rect 22714 82100 22733 82156
rect 22789 82100 22808 82156
rect 22714 82076 22808 82100
rect 22714 82020 22733 82076
rect 22789 82020 22808 82076
rect 22714 81996 22808 82020
rect 22714 81940 22733 81996
rect 22789 81940 22808 81996
rect 22714 81912 22808 81940
rect 25604 82236 25698 82264
rect 25604 82180 25623 82236
rect 25679 82180 25698 82236
rect 25604 82156 25698 82180
rect 25604 82100 25623 82156
rect 25679 82100 25698 82156
rect 25604 82076 25698 82100
rect 25604 82020 25623 82076
rect 25679 82020 25698 82076
rect 25604 81996 25698 82020
rect 25604 81940 25623 81996
rect 25679 81940 25698 81996
rect 25604 81912 25698 81940
rect 28494 82236 28588 82264
rect 28494 82180 28513 82236
rect 28569 82180 28588 82236
rect 28494 82156 28588 82180
rect 28494 82100 28513 82156
rect 28569 82100 28588 82156
rect 28494 82076 28588 82100
rect 28494 82020 28513 82076
rect 28569 82020 28588 82076
rect 28494 81996 28588 82020
rect 28494 81940 28513 81996
rect 28569 81940 28588 81996
rect 28494 81912 28588 81940
rect 31384 82236 31478 82264
rect 31384 82180 31403 82236
rect 31459 82180 31478 82236
rect 31384 82156 31478 82180
rect 31384 82100 31403 82156
rect 31459 82100 31478 82156
rect 31384 82076 31478 82100
rect 31384 82020 31403 82076
rect 31459 82020 31478 82076
rect 31384 81996 31478 82020
rect 31384 81940 31403 81996
rect 31459 81940 31478 81996
rect 31384 81912 31478 81940
rect 34274 82236 34368 82264
rect 34274 82180 34293 82236
rect 34349 82180 34368 82236
rect 34274 82156 34368 82180
rect 34274 82100 34293 82156
rect 34349 82100 34368 82156
rect 34274 82076 34368 82100
rect 34274 82020 34293 82076
rect 34349 82020 34368 82076
rect 34274 81996 34368 82020
rect 34274 81940 34293 81996
rect 34349 81940 34368 81996
rect 34274 81912 34368 81940
rect 37164 82236 37258 82264
rect 37164 82180 37183 82236
rect 37239 82180 37258 82236
rect 37164 82156 37258 82180
rect 37164 82100 37183 82156
rect 37239 82100 37258 82156
rect 37164 82076 37258 82100
rect 37164 82020 37183 82076
rect 37239 82020 37258 82076
rect 37164 81996 37258 82020
rect 37164 81940 37183 81996
rect 37239 81940 37258 81996
rect 37164 81912 37258 81940
rect 40054 82236 40148 82264
rect 40054 82180 40073 82236
rect 40129 82180 40148 82236
rect 40054 82156 40148 82180
rect 40054 82100 40073 82156
rect 40129 82100 40148 82156
rect 40054 82076 40148 82100
rect 40054 82020 40073 82076
rect 40129 82020 40148 82076
rect 40054 81996 40148 82020
rect 40054 81940 40073 81996
rect 40129 81940 40148 81996
rect 40054 81912 40148 81940
rect 42944 82236 43038 82264
rect 42944 82180 42963 82236
rect 43019 82180 43038 82236
rect 42944 82156 43038 82180
rect 42944 82100 42963 82156
rect 43019 82100 43038 82156
rect 42944 82076 43038 82100
rect 42944 82020 42963 82076
rect 43019 82020 43038 82076
rect 42944 81996 43038 82020
rect 42944 81940 42963 81996
rect 43019 81940 43038 81996
rect 42944 81912 43038 81940
rect 45834 82236 45928 82264
rect 45834 82180 45853 82236
rect 45909 82180 45928 82236
rect 45834 82156 45928 82180
rect 45834 82100 45853 82156
rect 45909 82100 45928 82156
rect 45834 82076 45928 82100
rect 45834 82020 45853 82076
rect 45909 82020 45928 82076
rect 45834 81996 45928 82020
rect 45834 81940 45853 81996
rect 45909 81940 45928 81996
rect 45834 81912 45928 81940
rect 48781 82236 48875 82264
rect 48781 82180 48800 82236
rect 48856 82180 48875 82236
rect 48781 82156 48875 82180
rect 48781 82100 48800 82156
rect 48856 82100 48875 82156
rect 48781 82076 48875 82100
rect 48781 82020 48800 82076
rect 48856 82020 48875 82076
rect 48781 81996 48875 82020
rect 48781 81940 48800 81996
rect 48856 81940 48875 81996
rect 48781 81912 48875 81940
rect 49630 82236 49830 82264
rect 49630 82180 49662 82236
rect 49718 82180 49742 82236
rect 49798 82180 49830 82236
rect 49630 82156 49830 82180
rect 49630 82100 49662 82156
rect 49718 82100 49742 82156
rect 49798 82100 49830 82156
rect 49630 82076 49830 82100
rect 49630 82020 49662 82076
rect 49718 82020 49742 82076
rect 49798 82020 49830 82076
rect 49630 81996 49830 82020
rect 49630 81940 49662 81996
rect 49718 81940 49742 81996
rect 49798 81940 49830 81996
rect 49630 81912 49830 81940
rect 52920 82236 53048 82264
rect 52920 82180 52956 82236
rect 53012 82180 53048 82236
rect 52920 82156 53048 82180
rect 52920 82100 52956 82156
rect 53012 82100 53048 82156
rect 52920 82076 53048 82100
rect 52920 82020 52956 82076
rect 53012 82020 53048 82076
rect 52920 81996 53048 82020
rect 52920 81940 52956 81996
rect 53012 81940 53048 81996
rect 52920 81912 53048 81940
rect 53078 82236 53206 82264
rect 53078 82180 53114 82236
rect 53170 82180 53206 82236
rect 53078 82156 53206 82180
rect 53078 82100 53114 82156
rect 53170 82100 53206 82156
rect 53078 82076 53206 82100
rect 53078 82020 53114 82076
rect 53170 82020 53206 82076
rect 53078 81996 53206 82020
rect 53078 81940 53114 81996
rect 53170 81940 53206 81996
rect 53078 81912 53206 81940
rect 53434 82236 53562 82264
rect 53434 82180 53470 82236
rect 53526 82180 53562 82236
rect 53434 82156 53562 82180
rect 53434 82100 53470 82156
rect 53526 82100 53562 82156
rect 53434 82076 53562 82100
rect 53434 82020 53470 82076
rect 53526 82020 53562 82076
rect 53434 81996 53562 82020
rect 53434 81940 53470 81996
rect 53526 81940 53562 81996
rect 53434 81912 53562 81940
rect 54752 82236 54880 82264
rect 54752 82180 54788 82236
rect 54844 82180 54880 82236
rect 54752 82156 54880 82180
rect 54752 82100 54788 82156
rect 54844 82100 54880 82156
rect 54752 82076 54880 82100
rect 54752 82020 54788 82076
rect 54844 82020 54880 82076
rect 54752 81996 54880 82020
rect 54752 81940 54788 81996
rect 54844 81940 54880 81996
rect 54752 81912 54880 81940
rect 55345 82236 55473 82264
rect 55345 82180 55381 82236
rect 55437 82180 55473 82236
rect 55345 82156 55473 82180
rect 55345 82100 55381 82156
rect 55437 82100 55473 82156
rect 55345 82076 55473 82100
rect 55345 82020 55381 82076
rect 55437 82020 55473 82076
rect 55345 81996 55473 82020
rect 55345 81940 55381 81996
rect 55437 81940 55473 81996
rect 55345 81912 55473 81940
rect 56491 82236 56619 82264
rect 56491 82180 56527 82236
rect 56583 82180 56619 82236
rect 56491 82156 56619 82180
rect 56491 82100 56527 82156
rect 56583 82100 56619 82156
rect 56491 82076 56619 82100
rect 56491 82020 56527 82076
rect 56583 82020 56619 82076
rect 56491 81996 56619 82020
rect 56491 81940 56527 81996
rect 56583 81940 56619 81996
rect 56491 81912 56619 81940
rect 57941 82236 58121 82264
rect 57941 82180 57963 82236
rect 58019 82180 58043 82236
rect 58099 82180 58121 82236
rect 57941 82156 58121 82180
rect 57941 82100 57963 82156
rect 58019 82100 58043 82156
rect 58099 82100 58121 82156
rect 57941 82076 58121 82100
rect 57941 82020 57963 82076
rect 58019 82020 58043 82076
rect 58099 82020 58121 82076
rect 57941 81996 58121 82020
rect 57941 81940 57963 81996
rect 58019 81940 58043 81996
rect 58099 81940 58121 81996
rect 57941 81912 58121 81940
rect 59164 82236 59304 82264
rect 59164 82180 59206 82236
rect 59262 82180 59304 82236
rect 59164 82156 59304 82180
rect 59164 82100 59206 82156
rect 59262 82100 59304 82156
rect 59164 82076 59304 82100
rect 59164 82020 59206 82076
rect 59262 82020 59304 82076
rect 59164 81996 59304 82020
rect 59164 81940 59206 81996
rect 59262 81940 59304 81996
rect 59164 81912 59304 81940
rect 59334 82236 59450 82264
rect 59334 82180 59364 82236
rect 59420 82180 59450 82236
rect 59334 82156 59450 82180
rect 59334 82100 59364 82156
rect 59420 82100 59450 82156
rect 59334 82076 59450 82100
rect 59334 82020 59364 82076
rect 59420 82020 59450 82076
rect 59334 81996 59450 82020
rect 59334 81940 59364 81996
rect 59420 81940 59450 81996
rect 59334 81912 59450 81940
rect 59642 82236 59758 82264
rect 59642 82180 59672 82236
rect 59728 82180 59758 82236
rect 59642 82156 59758 82180
rect 59642 82100 59672 82156
rect 59728 82100 59758 82156
rect 59642 82076 59758 82100
rect 59642 82020 59672 82076
rect 59728 82020 59758 82076
rect 59642 81996 59758 82020
rect 59642 81940 59672 81996
rect 59728 81940 59758 81996
rect 59642 81912 59758 81940
rect 59788 82236 59904 82264
rect 59788 82180 59818 82236
rect 59874 82180 59904 82236
rect 59788 82156 59904 82180
rect 59788 82100 59818 82156
rect 59874 82100 59904 82156
rect 59788 82076 59904 82100
rect 59788 82020 59818 82076
rect 59874 82020 59904 82076
rect 59788 81996 59904 82020
rect 59788 81940 59818 81996
rect 59874 81940 59904 81996
rect 59788 81912 59904 81940
rect 59934 82236 60110 82264
rect 59934 82180 59954 82236
rect 60010 82180 60034 82236
rect 60090 82180 60110 82236
rect 59934 82156 60110 82180
rect 59934 82100 59954 82156
rect 60010 82100 60034 82156
rect 60090 82100 60110 82156
rect 59934 82076 60110 82100
rect 59934 82020 59954 82076
rect 60010 82020 60034 82076
rect 60090 82020 60110 82076
rect 59934 81996 60110 82020
rect 59934 81940 59954 81996
rect 60010 81940 60034 81996
rect 60090 81940 60110 81996
rect 59934 81912 60110 81940
rect 62307 82236 62481 82264
rect 62307 82180 62326 82236
rect 62382 82180 62406 82236
rect 62462 82180 62481 82236
rect 62307 82156 62481 82180
rect 62307 82100 62326 82156
rect 62382 82100 62406 82156
rect 62462 82100 62481 82156
rect 62307 82076 62481 82100
rect 62307 82020 62326 82076
rect 62382 82020 62406 82076
rect 62462 82020 62481 82076
rect 62307 81996 62481 82020
rect 62307 81940 62326 81996
rect 62382 81940 62406 81996
rect 62462 81940 62481 81996
rect 62307 81912 62481 81940
rect 64892 81802 64920 84186
rect 71836 83258 72188 84294
rect 71836 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 72188 83258
rect 66996 83156 67048 83162
rect 66996 83098 67048 83104
rect 64880 81796 64932 81802
rect 64880 81738 64932 81744
rect 64892 79898 64920 81738
rect 64880 79892 64932 79898
rect 64880 79834 64932 79840
rect 64892 77722 64920 79834
rect 66444 78736 66496 78742
rect 66444 78678 66496 78684
rect 64880 77716 64932 77722
rect 64880 77658 64932 77664
rect 64892 75206 64920 77658
rect 66260 76560 66312 76566
rect 66260 76502 66312 76508
rect 64880 75200 64932 75206
rect 64880 75142 64932 75148
rect 2020 74588 2124 74616
rect 2020 74532 2044 74588
rect 2100 74532 2124 74588
rect 2020 74508 2124 74532
rect 2020 74452 2044 74508
rect 2100 74452 2124 74508
rect 2020 74428 2124 74452
rect 2020 74372 2044 74428
rect 2100 74372 2124 74428
rect 2020 74348 2124 74372
rect 2020 74292 2044 74348
rect 2100 74292 2124 74348
rect 2020 74264 2124 74292
rect 5521 74588 5615 74616
rect 5521 74532 5540 74588
rect 5596 74532 5615 74588
rect 5521 74508 5615 74532
rect 5521 74452 5540 74508
rect 5596 74452 5615 74508
rect 5521 74428 5615 74452
rect 5521 74372 5540 74428
rect 5596 74372 5615 74428
rect 5521 74348 5615 74372
rect 5521 74292 5540 74348
rect 5596 74292 5615 74348
rect 5521 74264 5615 74292
rect 8411 74588 8505 74616
rect 8411 74532 8430 74588
rect 8486 74532 8505 74588
rect 8411 74508 8505 74532
rect 8411 74452 8430 74508
rect 8486 74452 8505 74508
rect 8411 74428 8505 74452
rect 8411 74372 8430 74428
rect 8486 74372 8505 74428
rect 8411 74348 8505 74372
rect 8411 74292 8430 74348
rect 8486 74292 8505 74348
rect 8411 74264 8505 74292
rect 11301 74588 11395 74616
rect 11301 74532 11320 74588
rect 11376 74532 11395 74588
rect 11301 74508 11395 74532
rect 11301 74452 11320 74508
rect 11376 74452 11395 74508
rect 11301 74428 11395 74452
rect 11301 74372 11320 74428
rect 11376 74372 11395 74428
rect 11301 74348 11395 74372
rect 11301 74292 11320 74348
rect 11376 74292 11395 74348
rect 11301 74264 11395 74292
rect 14191 74588 14285 74616
rect 14191 74532 14210 74588
rect 14266 74532 14285 74588
rect 14191 74508 14285 74532
rect 14191 74452 14210 74508
rect 14266 74452 14285 74508
rect 14191 74428 14285 74452
rect 14191 74372 14210 74428
rect 14266 74372 14285 74428
rect 14191 74348 14285 74372
rect 14191 74292 14210 74348
rect 14266 74292 14285 74348
rect 14191 74264 14285 74292
rect 17081 74588 17175 74616
rect 17081 74532 17100 74588
rect 17156 74532 17175 74588
rect 17081 74508 17175 74532
rect 17081 74452 17100 74508
rect 17156 74452 17175 74508
rect 17081 74428 17175 74452
rect 17081 74372 17100 74428
rect 17156 74372 17175 74428
rect 17081 74348 17175 74372
rect 17081 74292 17100 74348
rect 17156 74292 17175 74348
rect 17081 74264 17175 74292
rect 19971 74588 20065 74616
rect 19971 74532 19990 74588
rect 20046 74532 20065 74588
rect 19971 74508 20065 74532
rect 19971 74452 19990 74508
rect 20046 74452 20065 74508
rect 19971 74428 20065 74452
rect 19971 74372 19990 74428
rect 20046 74372 20065 74428
rect 19971 74348 20065 74372
rect 19971 74292 19990 74348
rect 20046 74292 20065 74348
rect 19971 74264 20065 74292
rect 22861 74588 22955 74616
rect 22861 74532 22880 74588
rect 22936 74532 22955 74588
rect 22861 74508 22955 74532
rect 22861 74452 22880 74508
rect 22936 74452 22955 74508
rect 22861 74428 22955 74452
rect 22861 74372 22880 74428
rect 22936 74372 22955 74428
rect 22861 74348 22955 74372
rect 22861 74292 22880 74348
rect 22936 74292 22955 74348
rect 22861 74264 22955 74292
rect 25751 74588 25845 74616
rect 25751 74532 25770 74588
rect 25826 74532 25845 74588
rect 25751 74508 25845 74532
rect 25751 74452 25770 74508
rect 25826 74452 25845 74508
rect 25751 74428 25845 74452
rect 25751 74372 25770 74428
rect 25826 74372 25845 74428
rect 25751 74348 25845 74372
rect 25751 74292 25770 74348
rect 25826 74292 25845 74348
rect 25751 74264 25845 74292
rect 28641 74588 28735 74616
rect 28641 74532 28660 74588
rect 28716 74532 28735 74588
rect 28641 74508 28735 74532
rect 28641 74452 28660 74508
rect 28716 74452 28735 74508
rect 28641 74428 28735 74452
rect 28641 74372 28660 74428
rect 28716 74372 28735 74428
rect 28641 74348 28735 74372
rect 28641 74292 28660 74348
rect 28716 74292 28735 74348
rect 28641 74264 28735 74292
rect 31531 74588 31625 74616
rect 31531 74532 31550 74588
rect 31606 74532 31625 74588
rect 31531 74508 31625 74532
rect 31531 74452 31550 74508
rect 31606 74452 31625 74508
rect 31531 74428 31625 74452
rect 31531 74372 31550 74428
rect 31606 74372 31625 74428
rect 31531 74348 31625 74372
rect 31531 74292 31550 74348
rect 31606 74292 31625 74348
rect 31531 74264 31625 74292
rect 34421 74588 34515 74616
rect 34421 74532 34440 74588
rect 34496 74532 34515 74588
rect 34421 74508 34515 74532
rect 34421 74452 34440 74508
rect 34496 74452 34515 74508
rect 34421 74428 34515 74452
rect 34421 74372 34440 74428
rect 34496 74372 34515 74428
rect 34421 74348 34515 74372
rect 34421 74292 34440 74348
rect 34496 74292 34515 74348
rect 34421 74264 34515 74292
rect 37311 74588 37405 74616
rect 37311 74532 37330 74588
rect 37386 74532 37405 74588
rect 37311 74508 37405 74532
rect 37311 74452 37330 74508
rect 37386 74452 37405 74508
rect 37311 74428 37405 74452
rect 37311 74372 37330 74428
rect 37386 74372 37405 74428
rect 37311 74348 37405 74372
rect 37311 74292 37330 74348
rect 37386 74292 37405 74348
rect 37311 74264 37405 74292
rect 40201 74588 40295 74616
rect 40201 74532 40220 74588
rect 40276 74532 40295 74588
rect 40201 74508 40295 74532
rect 40201 74452 40220 74508
rect 40276 74452 40295 74508
rect 40201 74428 40295 74452
rect 40201 74372 40220 74428
rect 40276 74372 40295 74428
rect 40201 74348 40295 74372
rect 40201 74292 40220 74348
rect 40276 74292 40295 74348
rect 40201 74264 40295 74292
rect 43091 74588 43185 74616
rect 43091 74532 43110 74588
rect 43166 74532 43185 74588
rect 43091 74508 43185 74532
rect 43091 74452 43110 74508
rect 43166 74452 43185 74508
rect 43091 74428 43185 74452
rect 43091 74372 43110 74428
rect 43166 74372 43185 74428
rect 43091 74348 43185 74372
rect 43091 74292 43110 74348
rect 43166 74292 43185 74348
rect 43091 74264 43185 74292
rect 45981 74588 46075 74616
rect 45981 74532 46000 74588
rect 46056 74532 46075 74588
rect 45981 74508 46075 74532
rect 45981 74452 46000 74508
rect 46056 74452 46075 74508
rect 45981 74428 46075 74452
rect 45981 74372 46000 74428
rect 46056 74372 46075 74428
rect 45981 74348 46075 74372
rect 45981 74292 46000 74348
rect 46056 74292 46075 74348
rect 45981 74264 46075 74292
rect 48989 74588 49083 74616
rect 48989 74532 49008 74588
rect 49064 74532 49083 74588
rect 48989 74508 49083 74532
rect 48989 74452 49008 74508
rect 49064 74452 49083 74508
rect 48989 74428 49083 74452
rect 48989 74372 49008 74428
rect 49064 74372 49083 74428
rect 48989 74348 49083 74372
rect 48989 74292 49008 74348
rect 49064 74292 49083 74348
rect 48989 74264 49083 74292
rect 52210 74588 52320 74616
rect 52210 74532 52237 74588
rect 52293 74532 52320 74588
rect 52210 74508 52320 74532
rect 52210 74452 52237 74508
rect 52293 74452 52320 74508
rect 52210 74428 52320 74452
rect 52210 74372 52237 74428
rect 52293 74372 52320 74428
rect 52210 74348 52320 74372
rect 52210 74292 52237 74348
rect 52293 74292 52320 74348
rect 52210 74264 52320 74292
rect 53602 74588 53730 74616
rect 53602 74532 53638 74588
rect 53694 74532 53730 74588
rect 53602 74508 53730 74532
rect 53602 74452 53638 74508
rect 53694 74452 53730 74508
rect 53602 74428 53730 74452
rect 53602 74372 53638 74428
rect 53694 74372 53730 74428
rect 53602 74348 53730 74372
rect 53602 74292 53638 74348
rect 53694 74292 53730 74348
rect 53602 74264 53730 74292
rect 53770 74588 53898 74616
rect 53770 74532 53806 74588
rect 53862 74532 53898 74588
rect 53770 74508 53898 74532
rect 53770 74452 53806 74508
rect 53862 74452 53898 74508
rect 53770 74428 53898 74452
rect 53770 74372 53806 74428
rect 53862 74372 53898 74428
rect 53770 74348 53898 74372
rect 53770 74292 53806 74348
rect 53862 74292 53898 74348
rect 53770 74264 53898 74292
rect 54514 74588 54642 74616
rect 54514 74532 54550 74588
rect 54606 74532 54642 74588
rect 54514 74508 54642 74532
rect 54514 74452 54550 74508
rect 54606 74452 54642 74508
rect 54514 74428 54642 74452
rect 54514 74372 54550 74428
rect 54606 74372 54642 74428
rect 54514 74348 54642 74372
rect 54514 74292 54550 74348
rect 54606 74292 54642 74348
rect 54514 74264 54642 74292
rect 54910 74588 55026 74616
rect 54910 74532 54940 74588
rect 54996 74532 55026 74588
rect 54910 74508 55026 74532
rect 54910 74452 54940 74508
rect 54996 74452 55026 74508
rect 54910 74428 55026 74452
rect 54910 74372 54940 74428
rect 54996 74372 55026 74428
rect 54910 74348 55026 74372
rect 54910 74292 54940 74348
rect 54996 74292 55026 74348
rect 54910 74264 55026 74292
rect 55620 74588 55748 74616
rect 55620 74532 55656 74588
rect 55712 74532 55748 74588
rect 55620 74508 55748 74532
rect 55620 74452 55656 74508
rect 55712 74452 55748 74508
rect 55620 74428 55748 74452
rect 55620 74372 55656 74428
rect 55712 74372 55748 74428
rect 55620 74348 55748 74372
rect 55620 74292 55656 74348
rect 55712 74292 55748 74348
rect 55620 74264 55748 74292
rect 56198 74588 56326 74616
rect 56198 74532 56234 74588
rect 56290 74532 56326 74588
rect 56198 74508 56326 74532
rect 56198 74452 56234 74508
rect 56290 74452 56326 74508
rect 56198 74428 56326 74452
rect 56198 74372 56234 74428
rect 56290 74372 56326 74428
rect 56198 74348 56326 74372
rect 56198 74292 56234 74348
rect 56290 74292 56326 74348
rect 56198 74264 56326 74292
rect 56649 74588 56765 74616
rect 56649 74532 56679 74588
rect 56735 74532 56765 74588
rect 56649 74508 56765 74532
rect 56649 74452 56679 74508
rect 56735 74452 56765 74508
rect 56649 74428 56765 74452
rect 56649 74372 56679 74428
rect 56735 74372 56765 74428
rect 56649 74348 56765 74372
rect 56649 74292 56679 74348
rect 56735 74292 56765 74348
rect 56649 74264 56765 74292
rect 56953 74588 57069 74616
rect 56953 74532 56983 74588
rect 57039 74532 57069 74588
rect 56953 74508 57069 74532
rect 56953 74452 56983 74508
rect 57039 74452 57069 74508
rect 56953 74428 57069 74452
rect 56953 74372 56983 74428
rect 57039 74372 57069 74428
rect 56953 74348 57069 74372
rect 56953 74292 56983 74348
rect 57039 74292 57069 74348
rect 56953 74264 57069 74292
rect 57795 74588 57911 74616
rect 57795 74532 57825 74588
rect 57881 74532 57911 74588
rect 57795 74508 57911 74532
rect 57795 74452 57825 74508
rect 57881 74452 57911 74508
rect 57795 74428 57911 74452
rect 57795 74372 57825 74428
rect 57881 74372 57911 74428
rect 57795 74348 57911 74372
rect 57795 74292 57825 74348
rect 57881 74292 57911 74348
rect 57795 74264 57911 74292
rect 58461 74588 58525 74616
rect 58461 74532 58465 74588
rect 58521 74532 58525 74588
rect 58461 74508 58525 74532
rect 58461 74452 58465 74508
rect 58521 74452 58525 74508
rect 58461 74428 58525 74452
rect 58461 74372 58465 74428
rect 58521 74372 58525 74428
rect 58461 74348 58525 74372
rect 58461 74292 58465 74348
rect 58521 74292 58525 74348
rect 58461 74264 58525 74292
rect 59018 74588 59134 74616
rect 59018 74532 59048 74588
rect 59104 74532 59134 74588
rect 59018 74508 59134 74532
rect 59018 74452 59048 74508
rect 59104 74452 59134 74508
rect 59018 74428 59134 74452
rect 59018 74372 59048 74428
rect 59104 74372 59134 74428
rect 59018 74348 59134 74372
rect 59018 74292 59048 74348
rect 59104 74292 59134 74348
rect 59018 74264 59134 74292
rect 60296 74588 60412 74616
rect 60296 74532 60326 74588
rect 60382 74532 60412 74588
rect 60296 74508 60412 74532
rect 60296 74452 60326 74508
rect 60382 74452 60412 74508
rect 60296 74428 60412 74452
rect 60296 74372 60326 74428
rect 60382 74372 60412 74428
rect 60296 74348 60412 74372
rect 60296 74292 60326 74348
rect 60382 74292 60412 74348
rect 60296 74264 60412 74292
rect 60454 74588 60570 74616
rect 60454 74532 60484 74588
rect 60540 74532 60570 74588
rect 60454 74508 60570 74532
rect 60454 74452 60484 74508
rect 60540 74452 60570 74508
rect 60454 74428 60570 74452
rect 60454 74372 60484 74428
rect 60540 74372 60570 74428
rect 60454 74348 60570 74372
rect 60454 74292 60484 74348
rect 60540 74292 60570 74348
rect 60454 74264 60570 74292
rect 62509 74588 62683 74616
rect 62509 74532 62528 74588
rect 62584 74532 62608 74588
rect 62664 74532 62683 74588
rect 62509 74508 62683 74532
rect 62509 74452 62528 74508
rect 62584 74452 62608 74508
rect 62664 74452 62683 74508
rect 62509 74428 62683 74452
rect 62509 74372 62528 74428
rect 62584 74372 62608 74428
rect 62664 74372 62683 74428
rect 62509 74348 62683 74372
rect 62509 74292 62528 74348
rect 62584 74292 62608 74348
rect 62664 74292 62683 74348
rect 62509 74264 62683 74292
rect 64892 73234 64920 75142
rect 66168 74112 66220 74118
rect 66168 74054 66220 74060
rect 64880 73228 64932 73234
rect 64880 73170 64932 73176
rect 2152 72236 2352 72264
rect 2152 72180 2184 72236
rect 2240 72180 2264 72236
rect 2320 72180 2352 72236
rect 2152 72156 2352 72180
rect 2152 72100 2184 72156
rect 2240 72100 2264 72156
rect 2320 72100 2352 72156
rect 2152 72076 2352 72100
rect 2152 72020 2184 72076
rect 2240 72020 2264 72076
rect 2320 72020 2352 72076
rect 2152 71996 2352 72020
rect 2152 71940 2184 71996
rect 2240 71940 2264 71996
rect 2320 71940 2352 71996
rect 2152 71912 2352 71940
rect 5374 72236 5468 72264
rect 5374 72180 5393 72236
rect 5449 72180 5468 72236
rect 5374 72156 5468 72180
rect 5374 72100 5393 72156
rect 5449 72100 5468 72156
rect 5374 72076 5468 72100
rect 5374 72020 5393 72076
rect 5449 72020 5468 72076
rect 5374 71996 5468 72020
rect 5374 71940 5393 71996
rect 5449 71940 5468 71996
rect 5374 71912 5468 71940
rect 8264 72236 8358 72264
rect 8264 72180 8283 72236
rect 8339 72180 8358 72236
rect 8264 72156 8358 72180
rect 8264 72100 8283 72156
rect 8339 72100 8358 72156
rect 8264 72076 8358 72100
rect 8264 72020 8283 72076
rect 8339 72020 8358 72076
rect 8264 71996 8358 72020
rect 8264 71940 8283 71996
rect 8339 71940 8358 71996
rect 8264 71912 8358 71940
rect 11154 72236 11248 72264
rect 11154 72180 11173 72236
rect 11229 72180 11248 72236
rect 11154 72156 11248 72180
rect 11154 72100 11173 72156
rect 11229 72100 11248 72156
rect 11154 72076 11248 72100
rect 11154 72020 11173 72076
rect 11229 72020 11248 72076
rect 11154 71996 11248 72020
rect 11154 71940 11173 71996
rect 11229 71940 11248 71996
rect 11154 71912 11248 71940
rect 14044 72236 14138 72264
rect 14044 72180 14063 72236
rect 14119 72180 14138 72236
rect 14044 72156 14138 72180
rect 14044 72100 14063 72156
rect 14119 72100 14138 72156
rect 14044 72076 14138 72100
rect 14044 72020 14063 72076
rect 14119 72020 14138 72076
rect 14044 71996 14138 72020
rect 14044 71940 14063 71996
rect 14119 71940 14138 71996
rect 14044 71912 14138 71940
rect 16934 72236 17028 72264
rect 16934 72180 16953 72236
rect 17009 72180 17028 72236
rect 16934 72156 17028 72180
rect 16934 72100 16953 72156
rect 17009 72100 17028 72156
rect 16934 72076 17028 72100
rect 16934 72020 16953 72076
rect 17009 72020 17028 72076
rect 16934 71996 17028 72020
rect 16934 71940 16953 71996
rect 17009 71940 17028 71996
rect 16934 71912 17028 71940
rect 19824 72236 19918 72264
rect 19824 72180 19843 72236
rect 19899 72180 19918 72236
rect 19824 72156 19918 72180
rect 19824 72100 19843 72156
rect 19899 72100 19918 72156
rect 19824 72076 19918 72100
rect 19824 72020 19843 72076
rect 19899 72020 19918 72076
rect 19824 71996 19918 72020
rect 19824 71940 19843 71996
rect 19899 71940 19918 71996
rect 19824 71912 19918 71940
rect 22714 72236 22808 72264
rect 22714 72180 22733 72236
rect 22789 72180 22808 72236
rect 22714 72156 22808 72180
rect 22714 72100 22733 72156
rect 22789 72100 22808 72156
rect 22714 72076 22808 72100
rect 22714 72020 22733 72076
rect 22789 72020 22808 72076
rect 22714 71996 22808 72020
rect 22714 71940 22733 71996
rect 22789 71940 22808 71996
rect 22714 71912 22808 71940
rect 25604 72236 25698 72264
rect 25604 72180 25623 72236
rect 25679 72180 25698 72236
rect 25604 72156 25698 72180
rect 25604 72100 25623 72156
rect 25679 72100 25698 72156
rect 25604 72076 25698 72100
rect 25604 72020 25623 72076
rect 25679 72020 25698 72076
rect 25604 71996 25698 72020
rect 25604 71940 25623 71996
rect 25679 71940 25698 71996
rect 25604 71912 25698 71940
rect 28494 72236 28588 72264
rect 28494 72180 28513 72236
rect 28569 72180 28588 72236
rect 28494 72156 28588 72180
rect 28494 72100 28513 72156
rect 28569 72100 28588 72156
rect 28494 72076 28588 72100
rect 28494 72020 28513 72076
rect 28569 72020 28588 72076
rect 28494 71996 28588 72020
rect 28494 71940 28513 71996
rect 28569 71940 28588 71996
rect 28494 71912 28588 71940
rect 31384 72236 31478 72264
rect 31384 72180 31403 72236
rect 31459 72180 31478 72236
rect 31384 72156 31478 72180
rect 31384 72100 31403 72156
rect 31459 72100 31478 72156
rect 31384 72076 31478 72100
rect 31384 72020 31403 72076
rect 31459 72020 31478 72076
rect 31384 71996 31478 72020
rect 31384 71940 31403 71996
rect 31459 71940 31478 71996
rect 31384 71912 31478 71940
rect 34274 72236 34368 72264
rect 34274 72180 34293 72236
rect 34349 72180 34368 72236
rect 34274 72156 34368 72180
rect 34274 72100 34293 72156
rect 34349 72100 34368 72156
rect 34274 72076 34368 72100
rect 34274 72020 34293 72076
rect 34349 72020 34368 72076
rect 34274 71996 34368 72020
rect 34274 71940 34293 71996
rect 34349 71940 34368 71996
rect 34274 71912 34368 71940
rect 37164 72236 37258 72264
rect 37164 72180 37183 72236
rect 37239 72180 37258 72236
rect 37164 72156 37258 72180
rect 37164 72100 37183 72156
rect 37239 72100 37258 72156
rect 37164 72076 37258 72100
rect 37164 72020 37183 72076
rect 37239 72020 37258 72076
rect 37164 71996 37258 72020
rect 37164 71940 37183 71996
rect 37239 71940 37258 71996
rect 37164 71912 37258 71940
rect 40054 72236 40148 72264
rect 40054 72180 40073 72236
rect 40129 72180 40148 72236
rect 40054 72156 40148 72180
rect 40054 72100 40073 72156
rect 40129 72100 40148 72156
rect 40054 72076 40148 72100
rect 40054 72020 40073 72076
rect 40129 72020 40148 72076
rect 40054 71996 40148 72020
rect 40054 71940 40073 71996
rect 40129 71940 40148 71996
rect 40054 71912 40148 71940
rect 42944 72236 43038 72264
rect 42944 72180 42963 72236
rect 43019 72180 43038 72236
rect 42944 72156 43038 72180
rect 42944 72100 42963 72156
rect 43019 72100 43038 72156
rect 42944 72076 43038 72100
rect 42944 72020 42963 72076
rect 43019 72020 43038 72076
rect 42944 71996 43038 72020
rect 42944 71940 42963 71996
rect 43019 71940 43038 71996
rect 42944 71912 43038 71940
rect 45834 72236 45928 72264
rect 45834 72180 45853 72236
rect 45909 72180 45928 72236
rect 45834 72156 45928 72180
rect 45834 72100 45853 72156
rect 45909 72100 45928 72156
rect 45834 72076 45928 72100
rect 45834 72020 45853 72076
rect 45909 72020 45928 72076
rect 45834 71996 45928 72020
rect 45834 71940 45853 71996
rect 45909 71940 45928 71996
rect 45834 71912 45928 71940
rect 48781 72236 48875 72264
rect 48781 72180 48800 72236
rect 48856 72180 48875 72236
rect 48781 72156 48875 72180
rect 48781 72100 48800 72156
rect 48856 72100 48875 72156
rect 48781 72076 48875 72100
rect 48781 72020 48800 72076
rect 48856 72020 48875 72076
rect 48781 71996 48875 72020
rect 48781 71940 48800 71996
rect 48856 71940 48875 71996
rect 48781 71912 48875 71940
rect 49630 72236 49830 72264
rect 49630 72180 49662 72236
rect 49718 72180 49742 72236
rect 49798 72180 49830 72236
rect 49630 72156 49830 72180
rect 49630 72100 49662 72156
rect 49718 72100 49742 72156
rect 49798 72100 49830 72156
rect 49630 72076 49830 72100
rect 49630 72020 49662 72076
rect 49718 72020 49742 72076
rect 49798 72020 49830 72076
rect 49630 71996 49830 72020
rect 49630 71940 49662 71996
rect 49718 71940 49742 71996
rect 49798 71940 49830 71996
rect 49630 71912 49830 71940
rect 52920 72236 53048 72264
rect 52920 72180 52956 72236
rect 53012 72180 53048 72236
rect 52920 72156 53048 72180
rect 52920 72100 52956 72156
rect 53012 72100 53048 72156
rect 52920 72076 53048 72100
rect 52920 72020 52956 72076
rect 53012 72020 53048 72076
rect 52920 71996 53048 72020
rect 52920 71940 52956 71996
rect 53012 71940 53048 71996
rect 52920 71912 53048 71940
rect 53078 72236 53206 72264
rect 53078 72180 53114 72236
rect 53170 72180 53206 72236
rect 53078 72156 53206 72180
rect 53078 72100 53114 72156
rect 53170 72100 53206 72156
rect 53078 72076 53206 72100
rect 53078 72020 53114 72076
rect 53170 72020 53206 72076
rect 53078 71996 53206 72020
rect 53078 71940 53114 71996
rect 53170 71940 53206 71996
rect 53078 71912 53206 71940
rect 53434 72236 53562 72264
rect 53434 72180 53470 72236
rect 53526 72180 53562 72236
rect 53434 72156 53562 72180
rect 53434 72100 53470 72156
rect 53526 72100 53562 72156
rect 53434 72076 53562 72100
rect 53434 72020 53470 72076
rect 53526 72020 53562 72076
rect 53434 71996 53562 72020
rect 53434 71940 53470 71996
rect 53526 71940 53562 71996
rect 53434 71912 53562 71940
rect 54752 72236 54880 72264
rect 54752 72180 54788 72236
rect 54844 72180 54880 72236
rect 54752 72156 54880 72180
rect 54752 72100 54788 72156
rect 54844 72100 54880 72156
rect 54752 72076 54880 72100
rect 54752 72020 54788 72076
rect 54844 72020 54880 72076
rect 54752 71996 54880 72020
rect 54752 71940 54788 71996
rect 54844 71940 54880 71996
rect 54752 71912 54880 71940
rect 55345 72236 55473 72264
rect 55345 72180 55381 72236
rect 55437 72180 55473 72236
rect 55345 72156 55473 72180
rect 55345 72100 55381 72156
rect 55437 72100 55473 72156
rect 55345 72076 55473 72100
rect 55345 72020 55381 72076
rect 55437 72020 55473 72076
rect 55345 71996 55473 72020
rect 55345 71940 55381 71996
rect 55437 71940 55473 71996
rect 55345 71912 55473 71940
rect 56491 72236 56619 72264
rect 56491 72180 56527 72236
rect 56583 72180 56619 72236
rect 56491 72156 56619 72180
rect 56491 72100 56527 72156
rect 56583 72100 56619 72156
rect 56491 72076 56619 72100
rect 56491 72020 56527 72076
rect 56583 72020 56619 72076
rect 56491 71996 56619 72020
rect 56491 71940 56527 71996
rect 56583 71940 56619 71996
rect 56491 71912 56619 71940
rect 57941 72236 58121 72264
rect 57941 72180 57963 72236
rect 58019 72180 58043 72236
rect 58099 72180 58121 72236
rect 57941 72156 58121 72180
rect 57941 72100 57963 72156
rect 58019 72100 58043 72156
rect 58099 72100 58121 72156
rect 57941 72076 58121 72100
rect 57941 72020 57963 72076
rect 58019 72020 58043 72076
rect 58099 72020 58121 72076
rect 57941 71996 58121 72020
rect 57941 71940 57963 71996
rect 58019 71940 58043 71996
rect 58099 71940 58121 71996
rect 57941 71912 58121 71940
rect 59164 72236 59304 72264
rect 59164 72180 59206 72236
rect 59262 72180 59304 72236
rect 59164 72156 59304 72180
rect 59164 72100 59206 72156
rect 59262 72100 59304 72156
rect 59164 72076 59304 72100
rect 59164 72020 59206 72076
rect 59262 72020 59304 72076
rect 59164 71996 59304 72020
rect 59164 71940 59206 71996
rect 59262 71940 59304 71996
rect 59164 71912 59304 71940
rect 59334 72236 59450 72264
rect 59334 72180 59364 72236
rect 59420 72180 59450 72236
rect 59334 72156 59450 72180
rect 59334 72100 59364 72156
rect 59420 72100 59450 72156
rect 59334 72076 59450 72100
rect 59334 72020 59364 72076
rect 59420 72020 59450 72076
rect 59334 71996 59450 72020
rect 59334 71940 59364 71996
rect 59420 71940 59450 71996
rect 59334 71912 59450 71940
rect 59642 72236 59758 72264
rect 59642 72180 59672 72236
rect 59728 72180 59758 72236
rect 59642 72156 59758 72180
rect 59642 72100 59672 72156
rect 59728 72100 59758 72156
rect 59642 72076 59758 72100
rect 59642 72020 59672 72076
rect 59728 72020 59758 72076
rect 59642 71996 59758 72020
rect 59642 71940 59672 71996
rect 59728 71940 59758 71996
rect 59642 71912 59758 71940
rect 59788 72236 59904 72264
rect 59788 72180 59818 72236
rect 59874 72180 59904 72236
rect 59788 72156 59904 72180
rect 59788 72100 59818 72156
rect 59874 72100 59904 72156
rect 59788 72076 59904 72100
rect 59788 72020 59818 72076
rect 59874 72020 59904 72076
rect 59788 71996 59904 72020
rect 59788 71940 59818 71996
rect 59874 71940 59904 71996
rect 59788 71912 59904 71940
rect 59934 72236 60110 72264
rect 59934 72180 59954 72236
rect 60010 72180 60034 72236
rect 60090 72180 60110 72236
rect 59934 72156 60110 72180
rect 59934 72100 59954 72156
rect 60010 72100 60034 72156
rect 60090 72100 60110 72156
rect 59934 72076 60110 72100
rect 59934 72020 59954 72076
rect 60010 72020 60034 72076
rect 60090 72020 60110 72076
rect 59934 71996 60110 72020
rect 59934 71940 59954 71996
rect 60010 71940 60034 71996
rect 60090 71940 60110 71996
rect 59934 71912 60110 71940
rect 62307 72236 62481 72264
rect 62307 72180 62326 72236
rect 62382 72180 62406 72236
rect 62462 72180 62481 72236
rect 62307 72156 62481 72180
rect 62307 72100 62326 72156
rect 62382 72100 62406 72156
rect 62462 72100 62481 72156
rect 62307 72076 62481 72100
rect 62307 72020 62326 72076
rect 62382 72020 62406 72076
rect 62462 72020 62481 72076
rect 62307 71996 62481 72020
rect 62307 71940 62326 71996
rect 62382 71940 62406 71996
rect 62462 71940 62481 71996
rect 62307 71912 62481 71940
rect 64892 71126 64920 73170
rect 65064 71800 65116 71806
rect 65064 71742 65116 71748
rect 64880 71120 64932 71126
rect 64880 71062 64932 71068
rect 63684 69624 63736 69630
rect 63684 69566 63736 69572
rect 63500 67770 63552 67776
rect 63500 67712 63552 67718
rect 2020 64588 2124 64616
rect 2020 64532 2044 64588
rect 2100 64532 2124 64588
rect 2020 64508 2124 64532
rect 2020 64452 2044 64508
rect 2100 64452 2124 64508
rect 2020 64428 2124 64452
rect 2020 64372 2044 64428
rect 2100 64372 2124 64428
rect 2020 64348 2124 64372
rect 2020 64292 2044 64348
rect 2100 64292 2124 64348
rect 2020 64264 2124 64292
rect 5521 64588 5615 64616
rect 5521 64532 5540 64588
rect 5596 64532 5615 64588
rect 5521 64508 5615 64532
rect 5521 64452 5540 64508
rect 5596 64452 5615 64508
rect 5521 64428 5615 64452
rect 5521 64372 5540 64428
rect 5596 64372 5615 64428
rect 5521 64348 5615 64372
rect 5521 64292 5540 64348
rect 5596 64292 5615 64348
rect 5521 64264 5615 64292
rect 8411 64588 8505 64616
rect 8411 64532 8430 64588
rect 8486 64532 8505 64588
rect 8411 64508 8505 64532
rect 8411 64452 8430 64508
rect 8486 64452 8505 64508
rect 8411 64428 8505 64452
rect 8411 64372 8430 64428
rect 8486 64372 8505 64428
rect 8411 64348 8505 64372
rect 8411 64292 8430 64348
rect 8486 64292 8505 64348
rect 8411 64264 8505 64292
rect 11301 64588 11395 64616
rect 11301 64532 11320 64588
rect 11376 64532 11395 64588
rect 11301 64508 11395 64532
rect 11301 64452 11320 64508
rect 11376 64452 11395 64508
rect 11301 64428 11395 64452
rect 11301 64372 11320 64428
rect 11376 64372 11395 64428
rect 11301 64348 11395 64372
rect 11301 64292 11320 64348
rect 11376 64292 11395 64348
rect 11301 64264 11395 64292
rect 14191 64588 14285 64616
rect 14191 64532 14210 64588
rect 14266 64532 14285 64588
rect 14191 64508 14285 64532
rect 14191 64452 14210 64508
rect 14266 64452 14285 64508
rect 14191 64428 14285 64452
rect 14191 64372 14210 64428
rect 14266 64372 14285 64428
rect 14191 64348 14285 64372
rect 14191 64292 14210 64348
rect 14266 64292 14285 64348
rect 14191 64264 14285 64292
rect 17081 64588 17175 64616
rect 17081 64532 17100 64588
rect 17156 64532 17175 64588
rect 17081 64508 17175 64532
rect 17081 64452 17100 64508
rect 17156 64452 17175 64508
rect 17081 64428 17175 64452
rect 17081 64372 17100 64428
rect 17156 64372 17175 64428
rect 17081 64348 17175 64372
rect 17081 64292 17100 64348
rect 17156 64292 17175 64348
rect 17081 64264 17175 64292
rect 19971 64588 20065 64616
rect 19971 64532 19990 64588
rect 20046 64532 20065 64588
rect 19971 64508 20065 64532
rect 19971 64452 19990 64508
rect 20046 64452 20065 64508
rect 19971 64428 20065 64452
rect 19971 64372 19990 64428
rect 20046 64372 20065 64428
rect 19971 64348 20065 64372
rect 19971 64292 19990 64348
rect 20046 64292 20065 64348
rect 19971 64264 20065 64292
rect 22861 64588 22955 64616
rect 22861 64532 22880 64588
rect 22936 64532 22955 64588
rect 22861 64508 22955 64532
rect 22861 64452 22880 64508
rect 22936 64452 22955 64508
rect 22861 64428 22955 64452
rect 22861 64372 22880 64428
rect 22936 64372 22955 64428
rect 22861 64348 22955 64372
rect 22861 64292 22880 64348
rect 22936 64292 22955 64348
rect 22861 64264 22955 64292
rect 25751 64588 25845 64616
rect 25751 64532 25770 64588
rect 25826 64532 25845 64588
rect 25751 64508 25845 64532
rect 25751 64452 25770 64508
rect 25826 64452 25845 64508
rect 25751 64428 25845 64452
rect 25751 64372 25770 64428
rect 25826 64372 25845 64428
rect 25751 64348 25845 64372
rect 25751 64292 25770 64348
rect 25826 64292 25845 64348
rect 25751 64264 25845 64292
rect 28641 64588 28735 64616
rect 28641 64532 28660 64588
rect 28716 64532 28735 64588
rect 28641 64508 28735 64532
rect 28641 64452 28660 64508
rect 28716 64452 28735 64508
rect 28641 64428 28735 64452
rect 28641 64372 28660 64428
rect 28716 64372 28735 64428
rect 28641 64348 28735 64372
rect 28641 64292 28660 64348
rect 28716 64292 28735 64348
rect 28641 64264 28735 64292
rect 31531 64588 31625 64616
rect 31531 64532 31550 64588
rect 31606 64532 31625 64588
rect 31531 64508 31625 64532
rect 31531 64452 31550 64508
rect 31606 64452 31625 64508
rect 31531 64428 31625 64452
rect 31531 64372 31550 64428
rect 31606 64372 31625 64428
rect 31531 64348 31625 64372
rect 31531 64292 31550 64348
rect 31606 64292 31625 64348
rect 31531 64264 31625 64292
rect 34421 64588 34515 64616
rect 34421 64532 34440 64588
rect 34496 64532 34515 64588
rect 34421 64508 34515 64532
rect 34421 64452 34440 64508
rect 34496 64452 34515 64508
rect 34421 64428 34515 64452
rect 34421 64372 34440 64428
rect 34496 64372 34515 64428
rect 34421 64348 34515 64372
rect 34421 64292 34440 64348
rect 34496 64292 34515 64348
rect 34421 64264 34515 64292
rect 37311 64588 37405 64616
rect 37311 64532 37330 64588
rect 37386 64532 37405 64588
rect 37311 64508 37405 64532
rect 37311 64452 37330 64508
rect 37386 64452 37405 64508
rect 37311 64428 37405 64452
rect 37311 64372 37330 64428
rect 37386 64372 37405 64428
rect 37311 64348 37405 64372
rect 37311 64292 37330 64348
rect 37386 64292 37405 64348
rect 37311 64264 37405 64292
rect 40201 64588 40295 64616
rect 40201 64532 40220 64588
rect 40276 64532 40295 64588
rect 40201 64508 40295 64532
rect 40201 64452 40220 64508
rect 40276 64452 40295 64508
rect 40201 64428 40295 64452
rect 40201 64372 40220 64428
rect 40276 64372 40295 64428
rect 40201 64348 40295 64372
rect 40201 64292 40220 64348
rect 40276 64292 40295 64348
rect 40201 64264 40295 64292
rect 43091 64588 43185 64616
rect 43091 64532 43110 64588
rect 43166 64532 43185 64588
rect 43091 64508 43185 64532
rect 43091 64452 43110 64508
rect 43166 64452 43185 64508
rect 43091 64428 43185 64452
rect 43091 64372 43110 64428
rect 43166 64372 43185 64428
rect 43091 64348 43185 64372
rect 43091 64292 43110 64348
rect 43166 64292 43185 64348
rect 43091 64264 43185 64292
rect 45981 64588 46075 64616
rect 45981 64532 46000 64588
rect 46056 64532 46075 64588
rect 45981 64508 46075 64532
rect 45981 64452 46000 64508
rect 46056 64452 46075 64508
rect 45981 64428 46075 64452
rect 45981 64372 46000 64428
rect 46056 64372 46075 64428
rect 45981 64348 46075 64372
rect 45981 64292 46000 64348
rect 46056 64292 46075 64348
rect 45981 64264 46075 64292
rect 48989 64588 49083 64616
rect 48989 64532 49008 64588
rect 49064 64532 49083 64588
rect 48989 64508 49083 64532
rect 48989 64452 49008 64508
rect 49064 64452 49083 64508
rect 48989 64428 49083 64452
rect 48989 64372 49008 64428
rect 49064 64372 49083 64428
rect 48989 64348 49083 64372
rect 48989 64292 49008 64348
rect 49064 64292 49083 64348
rect 48989 64264 49083 64292
rect 52210 64588 52320 64616
rect 52210 64532 52237 64588
rect 52293 64532 52320 64588
rect 52210 64508 52320 64532
rect 52210 64452 52237 64508
rect 52293 64452 52320 64508
rect 52210 64428 52320 64452
rect 52210 64372 52237 64428
rect 52293 64372 52320 64428
rect 52210 64348 52320 64372
rect 52210 64292 52237 64348
rect 52293 64292 52320 64348
rect 52210 64264 52320 64292
rect 53602 64588 53730 64616
rect 53602 64532 53638 64588
rect 53694 64532 53730 64588
rect 53602 64508 53730 64532
rect 53602 64452 53638 64508
rect 53694 64452 53730 64508
rect 53602 64428 53730 64452
rect 53602 64372 53638 64428
rect 53694 64372 53730 64428
rect 53602 64348 53730 64372
rect 53602 64292 53638 64348
rect 53694 64292 53730 64348
rect 53602 64264 53730 64292
rect 53770 64588 53898 64616
rect 53770 64532 53806 64588
rect 53862 64532 53898 64588
rect 53770 64508 53898 64532
rect 53770 64452 53806 64508
rect 53862 64452 53898 64508
rect 53770 64428 53898 64452
rect 53770 64372 53806 64428
rect 53862 64372 53898 64428
rect 53770 64348 53898 64372
rect 53770 64292 53806 64348
rect 53862 64292 53898 64348
rect 53770 64264 53898 64292
rect 54514 64588 54642 64616
rect 54514 64532 54550 64588
rect 54606 64532 54642 64588
rect 54514 64508 54642 64532
rect 54514 64452 54550 64508
rect 54606 64452 54642 64508
rect 54514 64428 54642 64452
rect 54514 64372 54550 64428
rect 54606 64372 54642 64428
rect 54514 64348 54642 64372
rect 54514 64292 54550 64348
rect 54606 64292 54642 64348
rect 54514 64264 54642 64292
rect 54910 64588 55026 64616
rect 54910 64532 54940 64588
rect 54996 64532 55026 64588
rect 54910 64508 55026 64532
rect 54910 64452 54940 64508
rect 54996 64452 55026 64508
rect 54910 64428 55026 64452
rect 54910 64372 54940 64428
rect 54996 64372 55026 64428
rect 54910 64348 55026 64372
rect 54910 64292 54940 64348
rect 54996 64292 55026 64348
rect 54910 64264 55026 64292
rect 55620 64588 55748 64616
rect 55620 64532 55656 64588
rect 55712 64532 55748 64588
rect 55620 64508 55748 64532
rect 55620 64452 55656 64508
rect 55712 64452 55748 64508
rect 55620 64428 55748 64452
rect 55620 64372 55656 64428
rect 55712 64372 55748 64428
rect 55620 64348 55748 64372
rect 55620 64292 55656 64348
rect 55712 64292 55748 64348
rect 55620 64264 55748 64292
rect 56198 64588 56326 64616
rect 56198 64532 56234 64588
rect 56290 64532 56326 64588
rect 56198 64508 56326 64532
rect 56198 64452 56234 64508
rect 56290 64452 56326 64508
rect 56198 64428 56326 64452
rect 56198 64372 56234 64428
rect 56290 64372 56326 64428
rect 56198 64348 56326 64372
rect 56198 64292 56234 64348
rect 56290 64292 56326 64348
rect 56198 64264 56326 64292
rect 56649 64588 56765 64616
rect 56649 64532 56679 64588
rect 56735 64532 56765 64588
rect 56649 64508 56765 64532
rect 56649 64452 56679 64508
rect 56735 64452 56765 64508
rect 56649 64428 56765 64452
rect 56649 64372 56679 64428
rect 56735 64372 56765 64428
rect 56649 64348 56765 64372
rect 56649 64292 56679 64348
rect 56735 64292 56765 64348
rect 56649 64264 56765 64292
rect 56953 64588 57069 64616
rect 56953 64532 56983 64588
rect 57039 64532 57069 64588
rect 56953 64508 57069 64532
rect 56953 64452 56983 64508
rect 57039 64452 57069 64508
rect 56953 64428 57069 64452
rect 56953 64372 56983 64428
rect 57039 64372 57069 64428
rect 56953 64348 57069 64372
rect 56953 64292 56983 64348
rect 57039 64292 57069 64348
rect 56953 64264 57069 64292
rect 57795 64588 57911 64616
rect 57795 64532 57825 64588
rect 57881 64532 57911 64588
rect 57795 64508 57911 64532
rect 57795 64452 57825 64508
rect 57881 64452 57911 64508
rect 57795 64428 57911 64452
rect 57795 64372 57825 64428
rect 57881 64372 57911 64428
rect 57795 64348 57911 64372
rect 57795 64292 57825 64348
rect 57881 64292 57911 64348
rect 57795 64264 57911 64292
rect 58461 64588 58525 64616
rect 58461 64532 58465 64588
rect 58521 64532 58525 64588
rect 58461 64508 58525 64532
rect 58461 64452 58465 64508
rect 58521 64452 58525 64508
rect 58461 64428 58525 64452
rect 58461 64372 58465 64428
rect 58521 64372 58525 64428
rect 58461 64348 58525 64372
rect 58461 64292 58465 64348
rect 58521 64292 58525 64348
rect 58461 64264 58525 64292
rect 59018 64588 59134 64616
rect 59018 64532 59048 64588
rect 59104 64532 59134 64588
rect 59018 64508 59134 64532
rect 59018 64452 59048 64508
rect 59104 64452 59134 64508
rect 59018 64428 59134 64452
rect 59018 64372 59048 64428
rect 59104 64372 59134 64428
rect 59018 64348 59134 64372
rect 59018 64292 59048 64348
rect 59104 64292 59134 64348
rect 59018 64264 59134 64292
rect 60296 64588 60412 64616
rect 60296 64532 60326 64588
rect 60382 64532 60412 64588
rect 60296 64508 60412 64532
rect 60296 64452 60326 64508
rect 60382 64452 60412 64508
rect 60296 64428 60412 64452
rect 60296 64372 60326 64428
rect 60382 64372 60412 64428
rect 60296 64348 60412 64372
rect 60296 64292 60326 64348
rect 60382 64292 60412 64348
rect 60296 64264 60412 64292
rect 60454 64588 60570 64616
rect 60454 64532 60484 64588
rect 60540 64532 60570 64588
rect 60454 64508 60570 64532
rect 60454 64452 60484 64508
rect 60540 64452 60570 64508
rect 60454 64428 60570 64452
rect 60454 64372 60484 64428
rect 60540 64372 60570 64428
rect 60454 64348 60570 64372
rect 60454 64292 60484 64348
rect 60540 64292 60570 64348
rect 60454 64264 60570 64292
rect 62509 64588 62683 64616
rect 62509 64532 62528 64588
rect 62584 64532 62608 64588
rect 62664 64532 62683 64588
rect 62509 64508 62683 64532
rect 62509 64452 62528 64508
rect 62584 64452 62608 64508
rect 62664 64452 62683 64508
rect 62509 64428 62683 64452
rect 62509 64372 62528 64428
rect 62584 64372 62608 64428
rect 62664 64372 62683 64428
rect 62509 64348 62683 64372
rect 62509 64292 62528 64348
rect 62584 64292 62608 64348
rect 62664 64292 62683 64348
rect 62509 64264 62683 64292
rect 2152 62236 2352 62264
rect 2152 62180 2184 62236
rect 2240 62180 2264 62236
rect 2320 62180 2352 62236
rect 2152 62156 2352 62180
rect 2152 62100 2184 62156
rect 2240 62100 2264 62156
rect 2320 62100 2352 62156
rect 2152 62076 2352 62100
rect 2152 62020 2184 62076
rect 2240 62020 2264 62076
rect 2320 62020 2352 62076
rect 2152 61996 2352 62020
rect 2152 61940 2184 61996
rect 2240 61940 2264 61996
rect 2320 61940 2352 61996
rect 2152 61912 2352 61940
rect 5374 62236 5468 62264
rect 5374 62180 5393 62236
rect 5449 62180 5468 62236
rect 5374 62156 5468 62180
rect 5374 62100 5393 62156
rect 5449 62100 5468 62156
rect 5374 62076 5468 62100
rect 5374 62020 5393 62076
rect 5449 62020 5468 62076
rect 5374 61996 5468 62020
rect 5374 61940 5393 61996
rect 5449 61940 5468 61996
rect 5374 61912 5468 61940
rect 8264 62236 8358 62264
rect 8264 62180 8283 62236
rect 8339 62180 8358 62236
rect 8264 62156 8358 62180
rect 8264 62100 8283 62156
rect 8339 62100 8358 62156
rect 8264 62076 8358 62100
rect 8264 62020 8283 62076
rect 8339 62020 8358 62076
rect 8264 61996 8358 62020
rect 8264 61940 8283 61996
rect 8339 61940 8358 61996
rect 8264 61912 8358 61940
rect 11154 62236 11248 62264
rect 11154 62180 11173 62236
rect 11229 62180 11248 62236
rect 11154 62156 11248 62180
rect 11154 62100 11173 62156
rect 11229 62100 11248 62156
rect 11154 62076 11248 62100
rect 11154 62020 11173 62076
rect 11229 62020 11248 62076
rect 11154 61996 11248 62020
rect 11154 61940 11173 61996
rect 11229 61940 11248 61996
rect 11154 61912 11248 61940
rect 14044 62236 14138 62264
rect 14044 62180 14063 62236
rect 14119 62180 14138 62236
rect 14044 62156 14138 62180
rect 14044 62100 14063 62156
rect 14119 62100 14138 62156
rect 14044 62076 14138 62100
rect 14044 62020 14063 62076
rect 14119 62020 14138 62076
rect 14044 61996 14138 62020
rect 14044 61940 14063 61996
rect 14119 61940 14138 61996
rect 14044 61912 14138 61940
rect 16934 62236 17028 62264
rect 16934 62180 16953 62236
rect 17009 62180 17028 62236
rect 16934 62156 17028 62180
rect 16934 62100 16953 62156
rect 17009 62100 17028 62156
rect 16934 62076 17028 62100
rect 16934 62020 16953 62076
rect 17009 62020 17028 62076
rect 16934 61996 17028 62020
rect 16934 61940 16953 61996
rect 17009 61940 17028 61996
rect 16934 61912 17028 61940
rect 19824 62236 19918 62264
rect 19824 62180 19843 62236
rect 19899 62180 19918 62236
rect 19824 62156 19918 62180
rect 19824 62100 19843 62156
rect 19899 62100 19918 62156
rect 19824 62076 19918 62100
rect 19824 62020 19843 62076
rect 19899 62020 19918 62076
rect 19824 61996 19918 62020
rect 19824 61940 19843 61996
rect 19899 61940 19918 61996
rect 19824 61912 19918 61940
rect 22714 62236 22808 62264
rect 22714 62180 22733 62236
rect 22789 62180 22808 62236
rect 22714 62156 22808 62180
rect 22714 62100 22733 62156
rect 22789 62100 22808 62156
rect 22714 62076 22808 62100
rect 22714 62020 22733 62076
rect 22789 62020 22808 62076
rect 22714 61996 22808 62020
rect 22714 61940 22733 61996
rect 22789 61940 22808 61996
rect 22714 61912 22808 61940
rect 25604 62236 25698 62264
rect 25604 62180 25623 62236
rect 25679 62180 25698 62236
rect 25604 62156 25698 62180
rect 25604 62100 25623 62156
rect 25679 62100 25698 62156
rect 25604 62076 25698 62100
rect 25604 62020 25623 62076
rect 25679 62020 25698 62076
rect 25604 61996 25698 62020
rect 25604 61940 25623 61996
rect 25679 61940 25698 61996
rect 25604 61912 25698 61940
rect 28494 62236 28588 62264
rect 28494 62180 28513 62236
rect 28569 62180 28588 62236
rect 28494 62156 28588 62180
rect 28494 62100 28513 62156
rect 28569 62100 28588 62156
rect 28494 62076 28588 62100
rect 28494 62020 28513 62076
rect 28569 62020 28588 62076
rect 28494 61996 28588 62020
rect 28494 61940 28513 61996
rect 28569 61940 28588 61996
rect 28494 61912 28588 61940
rect 31384 62236 31478 62264
rect 31384 62180 31403 62236
rect 31459 62180 31478 62236
rect 31384 62156 31478 62180
rect 31384 62100 31403 62156
rect 31459 62100 31478 62156
rect 31384 62076 31478 62100
rect 31384 62020 31403 62076
rect 31459 62020 31478 62076
rect 31384 61996 31478 62020
rect 31384 61940 31403 61996
rect 31459 61940 31478 61996
rect 31384 61912 31478 61940
rect 34274 62236 34368 62264
rect 34274 62180 34293 62236
rect 34349 62180 34368 62236
rect 34274 62156 34368 62180
rect 34274 62100 34293 62156
rect 34349 62100 34368 62156
rect 34274 62076 34368 62100
rect 34274 62020 34293 62076
rect 34349 62020 34368 62076
rect 34274 61996 34368 62020
rect 34274 61940 34293 61996
rect 34349 61940 34368 61996
rect 34274 61912 34368 61940
rect 37164 62236 37258 62264
rect 37164 62180 37183 62236
rect 37239 62180 37258 62236
rect 37164 62156 37258 62180
rect 37164 62100 37183 62156
rect 37239 62100 37258 62156
rect 37164 62076 37258 62100
rect 37164 62020 37183 62076
rect 37239 62020 37258 62076
rect 37164 61996 37258 62020
rect 37164 61940 37183 61996
rect 37239 61940 37258 61996
rect 37164 61912 37258 61940
rect 40054 62236 40148 62264
rect 40054 62180 40073 62236
rect 40129 62180 40148 62236
rect 40054 62156 40148 62180
rect 40054 62100 40073 62156
rect 40129 62100 40148 62156
rect 40054 62076 40148 62100
rect 40054 62020 40073 62076
rect 40129 62020 40148 62076
rect 40054 61996 40148 62020
rect 40054 61940 40073 61996
rect 40129 61940 40148 61996
rect 40054 61912 40148 61940
rect 42944 62236 43038 62264
rect 42944 62180 42963 62236
rect 43019 62180 43038 62236
rect 42944 62156 43038 62180
rect 42944 62100 42963 62156
rect 43019 62100 43038 62156
rect 42944 62076 43038 62100
rect 42944 62020 42963 62076
rect 43019 62020 43038 62076
rect 42944 61996 43038 62020
rect 42944 61940 42963 61996
rect 43019 61940 43038 61996
rect 42944 61912 43038 61940
rect 45834 62236 45928 62264
rect 45834 62180 45853 62236
rect 45909 62180 45928 62236
rect 45834 62156 45928 62180
rect 45834 62100 45853 62156
rect 45909 62100 45928 62156
rect 45834 62076 45928 62100
rect 45834 62020 45853 62076
rect 45909 62020 45928 62076
rect 45834 61996 45928 62020
rect 45834 61940 45853 61996
rect 45909 61940 45928 61996
rect 45834 61912 45928 61940
rect 48781 62236 48875 62264
rect 48781 62180 48800 62236
rect 48856 62180 48875 62236
rect 48781 62156 48875 62180
rect 48781 62100 48800 62156
rect 48856 62100 48875 62156
rect 48781 62076 48875 62100
rect 48781 62020 48800 62076
rect 48856 62020 48875 62076
rect 48781 61996 48875 62020
rect 48781 61940 48800 61996
rect 48856 61940 48875 61996
rect 48781 61912 48875 61940
rect 49630 62236 49830 62264
rect 49630 62180 49662 62236
rect 49718 62180 49742 62236
rect 49798 62180 49830 62236
rect 49630 62156 49830 62180
rect 49630 62100 49662 62156
rect 49718 62100 49742 62156
rect 49798 62100 49830 62156
rect 49630 62076 49830 62100
rect 49630 62020 49662 62076
rect 49718 62020 49742 62076
rect 49798 62020 49830 62076
rect 49630 61996 49830 62020
rect 49630 61940 49662 61996
rect 49718 61940 49742 61996
rect 49798 61940 49830 61996
rect 49630 61912 49830 61940
rect 52920 62236 53048 62264
rect 52920 62180 52956 62236
rect 53012 62180 53048 62236
rect 52920 62156 53048 62180
rect 52920 62100 52956 62156
rect 53012 62100 53048 62156
rect 52920 62076 53048 62100
rect 52920 62020 52956 62076
rect 53012 62020 53048 62076
rect 52920 61996 53048 62020
rect 52920 61940 52956 61996
rect 53012 61940 53048 61996
rect 52920 61912 53048 61940
rect 53078 62236 53206 62264
rect 53078 62180 53114 62236
rect 53170 62180 53206 62236
rect 53078 62156 53206 62180
rect 53078 62100 53114 62156
rect 53170 62100 53206 62156
rect 53078 62076 53206 62100
rect 53078 62020 53114 62076
rect 53170 62020 53206 62076
rect 53078 61996 53206 62020
rect 53078 61940 53114 61996
rect 53170 61940 53206 61996
rect 53078 61912 53206 61940
rect 53434 62236 53562 62264
rect 53434 62180 53470 62236
rect 53526 62180 53562 62236
rect 53434 62156 53562 62180
rect 53434 62100 53470 62156
rect 53526 62100 53562 62156
rect 53434 62076 53562 62100
rect 53434 62020 53470 62076
rect 53526 62020 53562 62076
rect 53434 61996 53562 62020
rect 53434 61940 53470 61996
rect 53526 61940 53562 61996
rect 53434 61912 53562 61940
rect 54752 62236 54880 62264
rect 54752 62180 54788 62236
rect 54844 62180 54880 62236
rect 54752 62156 54880 62180
rect 54752 62100 54788 62156
rect 54844 62100 54880 62156
rect 54752 62076 54880 62100
rect 54752 62020 54788 62076
rect 54844 62020 54880 62076
rect 54752 61996 54880 62020
rect 54752 61940 54788 61996
rect 54844 61940 54880 61996
rect 54752 61912 54880 61940
rect 55345 62236 55473 62264
rect 55345 62180 55381 62236
rect 55437 62180 55473 62236
rect 55345 62156 55473 62180
rect 55345 62100 55381 62156
rect 55437 62100 55473 62156
rect 55345 62076 55473 62100
rect 55345 62020 55381 62076
rect 55437 62020 55473 62076
rect 55345 61996 55473 62020
rect 55345 61940 55381 61996
rect 55437 61940 55473 61996
rect 55345 61912 55473 61940
rect 56491 62236 56619 62264
rect 56491 62180 56527 62236
rect 56583 62180 56619 62236
rect 56491 62156 56619 62180
rect 56491 62100 56527 62156
rect 56583 62100 56619 62156
rect 56491 62076 56619 62100
rect 56491 62020 56527 62076
rect 56583 62020 56619 62076
rect 56491 61996 56619 62020
rect 56491 61940 56527 61996
rect 56583 61940 56619 61996
rect 56491 61912 56619 61940
rect 57941 62236 58121 62264
rect 57941 62180 57963 62236
rect 58019 62180 58043 62236
rect 58099 62180 58121 62236
rect 57941 62156 58121 62180
rect 57941 62100 57963 62156
rect 58019 62100 58043 62156
rect 58099 62100 58121 62156
rect 57941 62076 58121 62100
rect 57941 62020 57963 62076
rect 58019 62020 58043 62076
rect 58099 62020 58121 62076
rect 57941 61996 58121 62020
rect 57941 61940 57963 61996
rect 58019 61940 58043 61996
rect 58099 61940 58121 61996
rect 57941 61912 58121 61940
rect 59164 62236 59304 62264
rect 59164 62180 59206 62236
rect 59262 62180 59304 62236
rect 59164 62156 59304 62180
rect 59164 62100 59206 62156
rect 59262 62100 59304 62156
rect 59164 62076 59304 62100
rect 59164 62020 59206 62076
rect 59262 62020 59304 62076
rect 59164 61996 59304 62020
rect 59164 61940 59206 61996
rect 59262 61940 59304 61996
rect 59164 61912 59304 61940
rect 59334 62236 59450 62264
rect 59334 62180 59364 62236
rect 59420 62180 59450 62236
rect 59334 62156 59450 62180
rect 59334 62100 59364 62156
rect 59420 62100 59450 62156
rect 59334 62076 59450 62100
rect 59334 62020 59364 62076
rect 59420 62020 59450 62076
rect 59334 61996 59450 62020
rect 59334 61940 59364 61996
rect 59420 61940 59450 61996
rect 59334 61912 59450 61940
rect 59642 62236 59758 62264
rect 59642 62180 59672 62236
rect 59728 62180 59758 62236
rect 59642 62156 59758 62180
rect 59642 62100 59672 62156
rect 59728 62100 59758 62156
rect 59642 62076 59758 62100
rect 59642 62020 59672 62076
rect 59728 62020 59758 62076
rect 59642 61996 59758 62020
rect 59642 61940 59672 61996
rect 59728 61940 59758 61996
rect 59642 61912 59758 61940
rect 59788 62236 59904 62264
rect 59788 62180 59818 62236
rect 59874 62180 59904 62236
rect 59788 62156 59904 62180
rect 59788 62100 59818 62156
rect 59874 62100 59904 62156
rect 59788 62076 59904 62100
rect 59788 62020 59818 62076
rect 59874 62020 59904 62076
rect 59788 61996 59904 62020
rect 59788 61940 59818 61996
rect 59874 61940 59904 61996
rect 59788 61912 59904 61940
rect 59934 62236 60110 62264
rect 59934 62180 59954 62236
rect 60010 62180 60034 62236
rect 60090 62180 60110 62236
rect 59934 62156 60110 62180
rect 59934 62100 59954 62156
rect 60010 62100 60034 62156
rect 60090 62100 60110 62156
rect 59934 62076 60110 62100
rect 59934 62020 59954 62076
rect 60010 62020 60034 62076
rect 60090 62020 60110 62076
rect 59934 61996 60110 62020
rect 59934 61940 59954 61996
rect 60010 61940 60034 61996
rect 60090 61940 60110 61996
rect 59934 61912 60110 61940
rect 62307 62236 62481 62264
rect 62307 62180 62326 62236
rect 62382 62180 62406 62236
rect 62462 62180 62481 62236
rect 62307 62156 62481 62180
rect 62307 62100 62326 62156
rect 62382 62100 62406 62156
rect 62462 62100 62481 62156
rect 62307 62076 62481 62100
rect 62307 62020 62326 62076
rect 62382 62020 62406 62076
rect 62462 62020 62481 62076
rect 62307 61996 62481 62020
rect 62307 61940 62326 61996
rect 62382 61940 62406 61996
rect 62462 61940 62481 61996
rect 62307 61912 62481 61940
rect 2020 54588 2124 54616
rect 2020 54532 2044 54588
rect 2100 54532 2124 54588
rect 2020 54508 2124 54532
rect 2020 54452 2044 54508
rect 2100 54452 2124 54508
rect 2020 54428 2124 54452
rect 2020 54372 2044 54428
rect 2100 54372 2124 54428
rect 2020 54348 2124 54372
rect 2020 54292 2044 54348
rect 2100 54292 2124 54348
rect 2020 54264 2124 54292
rect 5521 54588 5615 54616
rect 5521 54532 5540 54588
rect 5596 54532 5615 54588
rect 5521 54508 5615 54532
rect 5521 54452 5540 54508
rect 5596 54452 5615 54508
rect 5521 54428 5615 54452
rect 5521 54372 5540 54428
rect 5596 54372 5615 54428
rect 5521 54348 5615 54372
rect 5521 54292 5540 54348
rect 5596 54292 5615 54348
rect 5521 54264 5615 54292
rect 8411 54588 8505 54616
rect 8411 54532 8430 54588
rect 8486 54532 8505 54588
rect 8411 54508 8505 54532
rect 8411 54452 8430 54508
rect 8486 54452 8505 54508
rect 8411 54428 8505 54452
rect 8411 54372 8430 54428
rect 8486 54372 8505 54428
rect 8411 54348 8505 54372
rect 8411 54292 8430 54348
rect 8486 54292 8505 54348
rect 8411 54264 8505 54292
rect 11301 54588 11395 54616
rect 11301 54532 11320 54588
rect 11376 54532 11395 54588
rect 11301 54508 11395 54532
rect 11301 54452 11320 54508
rect 11376 54452 11395 54508
rect 11301 54428 11395 54452
rect 11301 54372 11320 54428
rect 11376 54372 11395 54428
rect 11301 54348 11395 54372
rect 11301 54292 11320 54348
rect 11376 54292 11395 54348
rect 11301 54264 11395 54292
rect 14191 54588 14285 54616
rect 14191 54532 14210 54588
rect 14266 54532 14285 54588
rect 14191 54508 14285 54532
rect 14191 54452 14210 54508
rect 14266 54452 14285 54508
rect 14191 54428 14285 54452
rect 14191 54372 14210 54428
rect 14266 54372 14285 54428
rect 14191 54348 14285 54372
rect 14191 54292 14210 54348
rect 14266 54292 14285 54348
rect 14191 54264 14285 54292
rect 17081 54588 17175 54616
rect 17081 54532 17100 54588
rect 17156 54532 17175 54588
rect 17081 54508 17175 54532
rect 17081 54452 17100 54508
rect 17156 54452 17175 54508
rect 17081 54428 17175 54452
rect 17081 54372 17100 54428
rect 17156 54372 17175 54428
rect 17081 54348 17175 54372
rect 17081 54292 17100 54348
rect 17156 54292 17175 54348
rect 17081 54264 17175 54292
rect 19971 54588 20065 54616
rect 19971 54532 19990 54588
rect 20046 54532 20065 54588
rect 19971 54508 20065 54532
rect 19971 54452 19990 54508
rect 20046 54452 20065 54508
rect 19971 54428 20065 54452
rect 19971 54372 19990 54428
rect 20046 54372 20065 54428
rect 19971 54348 20065 54372
rect 19971 54292 19990 54348
rect 20046 54292 20065 54348
rect 19971 54264 20065 54292
rect 22861 54588 22955 54616
rect 22861 54532 22880 54588
rect 22936 54532 22955 54588
rect 22861 54508 22955 54532
rect 22861 54452 22880 54508
rect 22936 54452 22955 54508
rect 22861 54428 22955 54452
rect 22861 54372 22880 54428
rect 22936 54372 22955 54428
rect 22861 54348 22955 54372
rect 22861 54292 22880 54348
rect 22936 54292 22955 54348
rect 22861 54264 22955 54292
rect 25751 54588 25845 54616
rect 25751 54532 25770 54588
rect 25826 54532 25845 54588
rect 25751 54508 25845 54532
rect 25751 54452 25770 54508
rect 25826 54452 25845 54508
rect 25751 54428 25845 54452
rect 25751 54372 25770 54428
rect 25826 54372 25845 54428
rect 25751 54348 25845 54372
rect 25751 54292 25770 54348
rect 25826 54292 25845 54348
rect 25751 54264 25845 54292
rect 28641 54588 28735 54616
rect 28641 54532 28660 54588
rect 28716 54532 28735 54588
rect 28641 54508 28735 54532
rect 28641 54452 28660 54508
rect 28716 54452 28735 54508
rect 28641 54428 28735 54452
rect 28641 54372 28660 54428
rect 28716 54372 28735 54428
rect 28641 54348 28735 54372
rect 28641 54292 28660 54348
rect 28716 54292 28735 54348
rect 28641 54264 28735 54292
rect 31531 54588 31625 54616
rect 31531 54532 31550 54588
rect 31606 54532 31625 54588
rect 31531 54508 31625 54532
rect 31531 54452 31550 54508
rect 31606 54452 31625 54508
rect 31531 54428 31625 54452
rect 31531 54372 31550 54428
rect 31606 54372 31625 54428
rect 31531 54348 31625 54372
rect 31531 54292 31550 54348
rect 31606 54292 31625 54348
rect 31531 54264 31625 54292
rect 34421 54588 34515 54616
rect 34421 54532 34440 54588
rect 34496 54532 34515 54588
rect 34421 54508 34515 54532
rect 34421 54452 34440 54508
rect 34496 54452 34515 54508
rect 34421 54428 34515 54452
rect 34421 54372 34440 54428
rect 34496 54372 34515 54428
rect 34421 54348 34515 54372
rect 34421 54292 34440 54348
rect 34496 54292 34515 54348
rect 34421 54264 34515 54292
rect 37311 54588 37405 54616
rect 37311 54532 37330 54588
rect 37386 54532 37405 54588
rect 37311 54508 37405 54532
rect 37311 54452 37330 54508
rect 37386 54452 37405 54508
rect 37311 54428 37405 54452
rect 37311 54372 37330 54428
rect 37386 54372 37405 54428
rect 37311 54348 37405 54372
rect 37311 54292 37330 54348
rect 37386 54292 37405 54348
rect 37311 54264 37405 54292
rect 40201 54588 40295 54616
rect 40201 54532 40220 54588
rect 40276 54532 40295 54588
rect 40201 54508 40295 54532
rect 40201 54452 40220 54508
rect 40276 54452 40295 54508
rect 40201 54428 40295 54452
rect 40201 54372 40220 54428
rect 40276 54372 40295 54428
rect 40201 54348 40295 54372
rect 40201 54292 40220 54348
rect 40276 54292 40295 54348
rect 40201 54264 40295 54292
rect 43091 54588 43185 54616
rect 43091 54532 43110 54588
rect 43166 54532 43185 54588
rect 43091 54508 43185 54532
rect 43091 54452 43110 54508
rect 43166 54452 43185 54508
rect 43091 54428 43185 54452
rect 43091 54372 43110 54428
rect 43166 54372 43185 54428
rect 43091 54348 43185 54372
rect 43091 54292 43110 54348
rect 43166 54292 43185 54348
rect 43091 54264 43185 54292
rect 45981 54588 46075 54616
rect 45981 54532 46000 54588
rect 46056 54532 46075 54588
rect 45981 54508 46075 54532
rect 45981 54452 46000 54508
rect 46056 54452 46075 54508
rect 45981 54428 46075 54452
rect 45981 54372 46000 54428
rect 46056 54372 46075 54428
rect 45981 54348 46075 54372
rect 45981 54292 46000 54348
rect 46056 54292 46075 54348
rect 45981 54264 46075 54292
rect 48989 54588 49083 54616
rect 48989 54532 49008 54588
rect 49064 54532 49083 54588
rect 48989 54508 49083 54532
rect 48989 54452 49008 54508
rect 49064 54452 49083 54508
rect 48989 54428 49083 54452
rect 48989 54372 49008 54428
rect 49064 54372 49083 54428
rect 48989 54348 49083 54372
rect 48989 54292 49008 54348
rect 49064 54292 49083 54348
rect 48989 54264 49083 54292
rect 52210 54588 52320 54616
rect 52210 54532 52237 54588
rect 52293 54532 52320 54588
rect 52210 54508 52320 54532
rect 52210 54452 52237 54508
rect 52293 54452 52320 54508
rect 52210 54428 52320 54452
rect 52210 54372 52237 54428
rect 52293 54372 52320 54428
rect 52210 54348 52320 54372
rect 52210 54292 52237 54348
rect 52293 54292 52320 54348
rect 52210 54264 52320 54292
rect 53602 54588 53730 54616
rect 53602 54532 53638 54588
rect 53694 54532 53730 54588
rect 53602 54508 53730 54532
rect 53602 54452 53638 54508
rect 53694 54452 53730 54508
rect 53602 54428 53730 54452
rect 53602 54372 53638 54428
rect 53694 54372 53730 54428
rect 53602 54348 53730 54372
rect 53602 54292 53638 54348
rect 53694 54292 53730 54348
rect 53602 54264 53730 54292
rect 53770 54588 53898 54616
rect 53770 54532 53806 54588
rect 53862 54532 53898 54588
rect 53770 54508 53898 54532
rect 53770 54452 53806 54508
rect 53862 54452 53898 54508
rect 53770 54428 53898 54452
rect 53770 54372 53806 54428
rect 53862 54372 53898 54428
rect 53770 54348 53898 54372
rect 53770 54292 53806 54348
rect 53862 54292 53898 54348
rect 53770 54264 53898 54292
rect 54514 54588 54642 54616
rect 54514 54532 54550 54588
rect 54606 54532 54642 54588
rect 54514 54508 54642 54532
rect 54514 54452 54550 54508
rect 54606 54452 54642 54508
rect 54514 54428 54642 54452
rect 54514 54372 54550 54428
rect 54606 54372 54642 54428
rect 54514 54348 54642 54372
rect 54514 54292 54550 54348
rect 54606 54292 54642 54348
rect 54514 54264 54642 54292
rect 54910 54588 55026 54616
rect 54910 54532 54940 54588
rect 54996 54532 55026 54588
rect 54910 54508 55026 54532
rect 54910 54452 54940 54508
rect 54996 54452 55026 54508
rect 54910 54428 55026 54452
rect 54910 54372 54940 54428
rect 54996 54372 55026 54428
rect 54910 54348 55026 54372
rect 54910 54292 54940 54348
rect 54996 54292 55026 54348
rect 54910 54264 55026 54292
rect 55620 54588 55748 54616
rect 55620 54532 55656 54588
rect 55712 54532 55748 54588
rect 55620 54508 55748 54532
rect 55620 54452 55656 54508
rect 55712 54452 55748 54508
rect 55620 54428 55748 54452
rect 55620 54372 55656 54428
rect 55712 54372 55748 54428
rect 55620 54348 55748 54372
rect 55620 54292 55656 54348
rect 55712 54292 55748 54348
rect 55620 54264 55748 54292
rect 56198 54588 56326 54616
rect 56198 54532 56234 54588
rect 56290 54532 56326 54588
rect 56198 54508 56326 54532
rect 56198 54452 56234 54508
rect 56290 54452 56326 54508
rect 56198 54428 56326 54452
rect 56198 54372 56234 54428
rect 56290 54372 56326 54428
rect 56198 54348 56326 54372
rect 56198 54292 56234 54348
rect 56290 54292 56326 54348
rect 56198 54264 56326 54292
rect 56649 54588 56765 54616
rect 56649 54532 56679 54588
rect 56735 54532 56765 54588
rect 56649 54508 56765 54532
rect 56649 54452 56679 54508
rect 56735 54452 56765 54508
rect 56649 54428 56765 54452
rect 56649 54372 56679 54428
rect 56735 54372 56765 54428
rect 56649 54348 56765 54372
rect 56649 54292 56679 54348
rect 56735 54292 56765 54348
rect 56649 54264 56765 54292
rect 56953 54588 57069 54616
rect 56953 54532 56983 54588
rect 57039 54532 57069 54588
rect 56953 54508 57069 54532
rect 56953 54452 56983 54508
rect 57039 54452 57069 54508
rect 56953 54428 57069 54452
rect 56953 54372 56983 54428
rect 57039 54372 57069 54428
rect 56953 54348 57069 54372
rect 56953 54292 56983 54348
rect 57039 54292 57069 54348
rect 56953 54264 57069 54292
rect 57795 54588 57911 54616
rect 57795 54532 57825 54588
rect 57881 54532 57911 54588
rect 57795 54508 57911 54532
rect 57795 54452 57825 54508
rect 57881 54452 57911 54508
rect 57795 54428 57911 54452
rect 57795 54372 57825 54428
rect 57881 54372 57911 54428
rect 57795 54348 57911 54372
rect 57795 54292 57825 54348
rect 57881 54292 57911 54348
rect 57795 54264 57911 54292
rect 58461 54588 58525 54616
rect 58461 54532 58465 54588
rect 58521 54532 58525 54588
rect 58461 54508 58525 54532
rect 58461 54452 58465 54508
rect 58521 54452 58525 54508
rect 58461 54428 58525 54452
rect 58461 54372 58465 54428
rect 58521 54372 58525 54428
rect 58461 54348 58525 54372
rect 58461 54292 58465 54348
rect 58521 54292 58525 54348
rect 58461 54264 58525 54292
rect 59018 54588 59134 54616
rect 59018 54532 59048 54588
rect 59104 54532 59134 54588
rect 59018 54508 59134 54532
rect 59018 54452 59048 54508
rect 59104 54452 59134 54508
rect 59018 54428 59134 54452
rect 59018 54372 59048 54428
rect 59104 54372 59134 54428
rect 59018 54348 59134 54372
rect 59018 54292 59048 54348
rect 59104 54292 59134 54348
rect 59018 54264 59134 54292
rect 60296 54588 60412 54616
rect 60296 54532 60326 54588
rect 60382 54532 60412 54588
rect 60296 54508 60412 54532
rect 60296 54452 60326 54508
rect 60382 54452 60412 54508
rect 60296 54428 60412 54452
rect 60296 54372 60326 54428
rect 60382 54372 60412 54428
rect 60296 54348 60412 54372
rect 60296 54292 60326 54348
rect 60382 54292 60412 54348
rect 60296 54264 60412 54292
rect 60454 54588 60570 54616
rect 60454 54532 60484 54588
rect 60540 54532 60570 54588
rect 60454 54508 60570 54532
rect 60454 54452 60484 54508
rect 60540 54452 60570 54508
rect 60454 54428 60570 54452
rect 60454 54372 60484 54428
rect 60540 54372 60570 54428
rect 60454 54348 60570 54372
rect 60454 54292 60484 54348
rect 60540 54292 60570 54348
rect 60454 54264 60570 54292
rect 62509 54588 62683 54616
rect 62509 54532 62528 54588
rect 62584 54532 62608 54588
rect 62664 54532 62683 54588
rect 62509 54508 62683 54532
rect 62509 54452 62528 54508
rect 62584 54452 62608 54508
rect 62664 54452 62683 54508
rect 62509 54428 62683 54452
rect 62509 54372 62528 54428
rect 62584 54372 62608 54428
rect 62664 54372 62683 54428
rect 62509 54348 62683 54372
rect 62509 54292 62528 54348
rect 62584 54292 62608 54348
rect 62664 54292 62683 54348
rect 62509 54264 62683 54292
rect 2152 52236 2352 52264
rect 2152 52180 2184 52236
rect 2240 52180 2264 52236
rect 2320 52180 2352 52236
rect 2152 52156 2352 52180
rect 2152 52100 2184 52156
rect 2240 52100 2264 52156
rect 2320 52100 2352 52156
rect 2152 52076 2352 52100
rect 2152 52020 2184 52076
rect 2240 52020 2264 52076
rect 2320 52020 2352 52076
rect 2152 51996 2352 52020
rect 2152 51940 2184 51996
rect 2240 51940 2264 51996
rect 2320 51940 2352 51996
rect 2152 51912 2352 51940
rect 5374 52236 5468 52264
rect 5374 52180 5393 52236
rect 5449 52180 5468 52236
rect 5374 52156 5468 52180
rect 5374 52100 5393 52156
rect 5449 52100 5468 52156
rect 5374 52076 5468 52100
rect 5374 52020 5393 52076
rect 5449 52020 5468 52076
rect 5374 51996 5468 52020
rect 5374 51940 5393 51996
rect 5449 51940 5468 51996
rect 5374 51912 5468 51940
rect 8264 52236 8358 52264
rect 8264 52180 8283 52236
rect 8339 52180 8358 52236
rect 8264 52156 8358 52180
rect 8264 52100 8283 52156
rect 8339 52100 8358 52156
rect 8264 52076 8358 52100
rect 8264 52020 8283 52076
rect 8339 52020 8358 52076
rect 8264 51996 8358 52020
rect 8264 51940 8283 51996
rect 8339 51940 8358 51996
rect 8264 51912 8358 51940
rect 11154 52236 11248 52264
rect 11154 52180 11173 52236
rect 11229 52180 11248 52236
rect 11154 52156 11248 52180
rect 11154 52100 11173 52156
rect 11229 52100 11248 52156
rect 11154 52076 11248 52100
rect 11154 52020 11173 52076
rect 11229 52020 11248 52076
rect 11154 51996 11248 52020
rect 11154 51940 11173 51996
rect 11229 51940 11248 51996
rect 11154 51912 11248 51940
rect 14044 52236 14138 52264
rect 14044 52180 14063 52236
rect 14119 52180 14138 52236
rect 14044 52156 14138 52180
rect 14044 52100 14063 52156
rect 14119 52100 14138 52156
rect 14044 52076 14138 52100
rect 14044 52020 14063 52076
rect 14119 52020 14138 52076
rect 14044 51996 14138 52020
rect 14044 51940 14063 51996
rect 14119 51940 14138 51996
rect 14044 51912 14138 51940
rect 16934 52236 17028 52264
rect 16934 52180 16953 52236
rect 17009 52180 17028 52236
rect 16934 52156 17028 52180
rect 16934 52100 16953 52156
rect 17009 52100 17028 52156
rect 16934 52076 17028 52100
rect 16934 52020 16953 52076
rect 17009 52020 17028 52076
rect 16934 51996 17028 52020
rect 16934 51940 16953 51996
rect 17009 51940 17028 51996
rect 16934 51912 17028 51940
rect 19824 52236 19918 52264
rect 19824 52180 19843 52236
rect 19899 52180 19918 52236
rect 19824 52156 19918 52180
rect 19824 52100 19843 52156
rect 19899 52100 19918 52156
rect 19824 52076 19918 52100
rect 19824 52020 19843 52076
rect 19899 52020 19918 52076
rect 19824 51996 19918 52020
rect 19824 51940 19843 51996
rect 19899 51940 19918 51996
rect 19824 51912 19918 51940
rect 22714 52236 22808 52264
rect 22714 52180 22733 52236
rect 22789 52180 22808 52236
rect 22714 52156 22808 52180
rect 22714 52100 22733 52156
rect 22789 52100 22808 52156
rect 22714 52076 22808 52100
rect 22714 52020 22733 52076
rect 22789 52020 22808 52076
rect 22714 51996 22808 52020
rect 22714 51940 22733 51996
rect 22789 51940 22808 51996
rect 22714 51912 22808 51940
rect 25604 52236 25698 52264
rect 25604 52180 25623 52236
rect 25679 52180 25698 52236
rect 25604 52156 25698 52180
rect 25604 52100 25623 52156
rect 25679 52100 25698 52156
rect 25604 52076 25698 52100
rect 25604 52020 25623 52076
rect 25679 52020 25698 52076
rect 25604 51996 25698 52020
rect 25604 51940 25623 51996
rect 25679 51940 25698 51996
rect 25604 51912 25698 51940
rect 28494 52236 28588 52264
rect 28494 52180 28513 52236
rect 28569 52180 28588 52236
rect 28494 52156 28588 52180
rect 28494 52100 28513 52156
rect 28569 52100 28588 52156
rect 28494 52076 28588 52100
rect 28494 52020 28513 52076
rect 28569 52020 28588 52076
rect 28494 51996 28588 52020
rect 28494 51940 28513 51996
rect 28569 51940 28588 51996
rect 28494 51912 28588 51940
rect 31384 52236 31478 52264
rect 31384 52180 31403 52236
rect 31459 52180 31478 52236
rect 31384 52156 31478 52180
rect 31384 52100 31403 52156
rect 31459 52100 31478 52156
rect 31384 52076 31478 52100
rect 31384 52020 31403 52076
rect 31459 52020 31478 52076
rect 31384 51996 31478 52020
rect 31384 51940 31403 51996
rect 31459 51940 31478 51996
rect 31384 51912 31478 51940
rect 34274 52236 34368 52264
rect 34274 52180 34293 52236
rect 34349 52180 34368 52236
rect 34274 52156 34368 52180
rect 34274 52100 34293 52156
rect 34349 52100 34368 52156
rect 34274 52076 34368 52100
rect 34274 52020 34293 52076
rect 34349 52020 34368 52076
rect 34274 51996 34368 52020
rect 34274 51940 34293 51996
rect 34349 51940 34368 51996
rect 34274 51912 34368 51940
rect 37164 52236 37258 52264
rect 37164 52180 37183 52236
rect 37239 52180 37258 52236
rect 37164 52156 37258 52180
rect 37164 52100 37183 52156
rect 37239 52100 37258 52156
rect 37164 52076 37258 52100
rect 37164 52020 37183 52076
rect 37239 52020 37258 52076
rect 37164 51996 37258 52020
rect 37164 51940 37183 51996
rect 37239 51940 37258 51996
rect 37164 51912 37258 51940
rect 40054 52236 40148 52264
rect 40054 52180 40073 52236
rect 40129 52180 40148 52236
rect 40054 52156 40148 52180
rect 40054 52100 40073 52156
rect 40129 52100 40148 52156
rect 40054 52076 40148 52100
rect 40054 52020 40073 52076
rect 40129 52020 40148 52076
rect 40054 51996 40148 52020
rect 40054 51940 40073 51996
rect 40129 51940 40148 51996
rect 40054 51912 40148 51940
rect 42944 52236 43038 52264
rect 42944 52180 42963 52236
rect 43019 52180 43038 52236
rect 42944 52156 43038 52180
rect 42944 52100 42963 52156
rect 43019 52100 43038 52156
rect 42944 52076 43038 52100
rect 42944 52020 42963 52076
rect 43019 52020 43038 52076
rect 42944 51996 43038 52020
rect 42944 51940 42963 51996
rect 43019 51940 43038 51996
rect 42944 51912 43038 51940
rect 45834 52236 45928 52264
rect 45834 52180 45853 52236
rect 45909 52180 45928 52236
rect 45834 52156 45928 52180
rect 45834 52100 45853 52156
rect 45909 52100 45928 52156
rect 45834 52076 45928 52100
rect 45834 52020 45853 52076
rect 45909 52020 45928 52076
rect 45834 51996 45928 52020
rect 45834 51940 45853 51996
rect 45909 51940 45928 51996
rect 45834 51912 45928 51940
rect 48781 52236 48875 52264
rect 48781 52180 48800 52236
rect 48856 52180 48875 52236
rect 48781 52156 48875 52180
rect 48781 52100 48800 52156
rect 48856 52100 48875 52156
rect 48781 52076 48875 52100
rect 48781 52020 48800 52076
rect 48856 52020 48875 52076
rect 48781 51996 48875 52020
rect 48781 51940 48800 51996
rect 48856 51940 48875 51996
rect 48781 51912 48875 51940
rect 49630 52236 49830 52264
rect 49630 52180 49662 52236
rect 49718 52180 49742 52236
rect 49798 52180 49830 52236
rect 49630 52156 49830 52180
rect 49630 52100 49662 52156
rect 49718 52100 49742 52156
rect 49798 52100 49830 52156
rect 49630 52076 49830 52100
rect 49630 52020 49662 52076
rect 49718 52020 49742 52076
rect 49798 52020 49830 52076
rect 49630 51996 49830 52020
rect 49630 51940 49662 51996
rect 49718 51940 49742 51996
rect 49798 51940 49830 51996
rect 49630 51912 49830 51940
rect 52920 52236 53048 52264
rect 52920 52180 52956 52236
rect 53012 52180 53048 52236
rect 52920 52156 53048 52180
rect 52920 52100 52956 52156
rect 53012 52100 53048 52156
rect 52920 52076 53048 52100
rect 52920 52020 52956 52076
rect 53012 52020 53048 52076
rect 52920 51996 53048 52020
rect 52920 51940 52956 51996
rect 53012 51940 53048 51996
rect 52920 51912 53048 51940
rect 53078 52236 53206 52264
rect 53078 52180 53114 52236
rect 53170 52180 53206 52236
rect 53078 52156 53206 52180
rect 53078 52100 53114 52156
rect 53170 52100 53206 52156
rect 53078 52076 53206 52100
rect 53078 52020 53114 52076
rect 53170 52020 53206 52076
rect 53078 51996 53206 52020
rect 53078 51940 53114 51996
rect 53170 51940 53206 51996
rect 53078 51912 53206 51940
rect 53434 52236 53562 52264
rect 53434 52180 53470 52236
rect 53526 52180 53562 52236
rect 53434 52156 53562 52180
rect 53434 52100 53470 52156
rect 53526 52100 53562 52156
rect 53434 52076 53562 52100
rect 53434 52020 53470 52076
rect 53526 52020 53562 52076
rect 53434 51996 53562 52020
rect 53434 51940 53470 51996
rect 53526 51940 53562 51996
rect 53434 51912 53562 51940
rect 54752 52236 54880 52264
rect 54752 52180 54788 52236
rect 54844 52180 54880 52236
rect 54752 52156 54880 52180
rect 54752 52100 54788 52156
rect 54844 52100 54880 52156
rect 54752 52076 54880 52100
rect 54752 52020 54788 52076
rect 54844 52020 54880 52076
rect 54752 51996 54880 52020
rect 54752 51940 54788 51996
rect 54844 51940 54880 51996
rect 54752 51912 54880 51940
rect 55345 52236 55473 52264
rect 55345 52180 55381 52236
rect 55437 52180 55473 52236
rect 55345 52156 55473 52180
rect 55345 52100 55381 52156
rect 55437 52100 55473 52156
rect 55345 52076 55473 52100
rect 55345 52020 55381 52076
rect 55437 52020 55473 52076
rect 55345 51996 55473 52020
rect 55345 51940 55381 51996
rect 55437 51940 55473 51996
rect 55345 51912 55473 51940
rect 56491 52236 56619 52264
rect 56491 52180 56527 52236
rect 56583 52180 56619 52236
rect 56491 52156 56619 52180
rect 56491 52100 56527 52156
rect 56583 52100 56619 52156
rect 56491 52076 56619 52100
rect 56491 52020 56527 52076
rect 56583 52020 56619 52076
rect 56491 51996 56619 52020
rect 56491 51940 56527 51996
rect 56583 51940 56619 51996
rect 56491 51912 56619 51940
rect 57941 52236 58121 52264
rect 57941 52180 57963 52236
rect 58019 52180 58043 52236
rect 58099 52180 58121 52236
rect 57941 52156 58121 52180
rect 57941 52100 57963 52156
rect 58019 52100 58043 52156
rect 58099 52100 58121 52156
rect 57941 52076 58121 52100
rect 57941 52020 57963 52076
rect 58019 52020 58043 52076
rect 58099 52020 58121 52076
rect 57941 51996 58121 52020
rect 57941 51940 57963 51996
rect 58019 51940 58043 51996
rect 58099 51940 58121 51996
rect 57941 51912 58121 51940
rect 59164 52236 59304 52264
rect 59164 52180 59206 52236
rect 59262 52180 59304 52236
rect 59164 52156 59304 52180
rect 59164 52100 59206 52156
rect 59262 52100 59304 52156
rect 59164 52076 59304 52100
rect 59164 52020 59206 52076
rect 59262 52020 59304 52076
rect 59164 51996 59304 52020
rect 59164 51940 59206 51996
rect 59262 51940 59304 51996
rect 59164 51912 59304 51940
rect 59334 52236 59450 52264
rect 59334 52180 59364 52236
rect 59420 52180 59450 52236
rect 59334 52156 59450 52180
rect 59334 52100 59364 52156
rect 59420 52100 59450 52156
rect 59334 52076 59450 52100
rect 59334 52020 59364 52076
rect 59420 52020 59450 52076
rect 59334 51996 59450 52020
rect 59334 51940 59364 51996
rect 59420 51940 59450 51996
rect 59334 51912 59450 51940
rect 59642 52236 59758 52264
rect 59642 52180 59672 52236
rect 59728 52180 59758 52236
rect 59642 52156 59758 52180
rect 59642 52100 59672 52156
rect 59728 52100 59758 52156
rect 59642 52076 59758 52100
rect 59642 52020 59672 52076
rect 59728 52020 59758 52076
rect 59642 51996 59758 52020
rect 59642 51940 59672 51996
rect 59728 51940 59758 51996
rect 59642 51912 59758 51940
rect 59788 52236 59904 52264
rect 59788 52180 59818 52236
rect 59874 52180 59904 52236
rect 59788 52156 59904 52180
rect 59788 52100 59818 52156
rect 59874 52100 59904 52156
rect 59788 52076 59904 52100
rect 59788 52020 59818 52076
rect 59874 52020 59904 52076
rect 59788 51996 59904 52020
rect 59788 51940 59818 51996
rect 59874 51940 59904 51996
rect 59788 51912 59904 51940
rect 59934 52236 60110 52264
rect 59934 52180 59954 52236
rect 60010 52180 60034 52236
rect 60090 52180 60110 52236
rect 59934 52156 60110 52180
rect 59934 52100 59954 52156
rect 60010 52100 60034 52156
rect 60090 52100 60110 52156
rect 59934 52076 60110 52100
rect 59934 52020 59954 52076
rect 60010 52020 60034 52076
rect 60090 52020 60110 52076
rect 59934 51996 60110 52020
rect 59934 51940 59954 51996
rect 60010 51940 60034 51996
rect 60090 51940 60110 51996
rect 59934 51912 60110 51940
rect 62307 52236 62481 52264
rect 62307 52180 62326 52236
rect 62382 52180 62406 52236
rect 62462 52180 62481 52236
rect 62307 52156 62481 52180
rect 62307 52100 62326 52156
rect 62382 52100 62406 52156
rect 62462 52100 62481 52156
rect 62307 52076 62481 52100
rect 62307 52020 62326 52076
rect 62382 52020 62406 52076
rect 62462 52020 62481 52076
rect 62307 51996 62481 52020
rect 62307 51940 62326 51996
rect 62382 51940 62406 51996
rect 62462 51940 62481 51996
rect 62307 51912 62481 51940
rect 2020 44588 2124 44616
rect 2020 44532 2044 44588
rect 2100 44532 2124 44588
rect 2020 44508 2124 44532
rect 2020 44452 2044 44508
rect 2100 44452 2124 44508
rect 2020 44428 2124 44452
rect 2020 44372 2044 44428
rect 2100 44372 2124 44428
rect 2020 44348 2124 44372
rect 2020 44292 2044 44348
rect 2100 44292 2124 44348
rect 2020 44264 2124 44292
rect 5521 44588 5615 44616
rect 5521 44532 5540 44588
rect 5596 44532 5615 44588
rect 5521 44508 5615 44532
rect 5521 44452 5540 44508
rect 5596 44452 5615 44508
rect 5521 44428 5615 44452
rect 5521 44372 5540 44428
rect 5596 44372 5615 44428
rect 5521 44348 5615 44372
rect 5521 44292 5540 44348
rect 5596 44292 5615 44348
rect 5521 44264 5615 44292
rect 8411 44588 8505 44616
rect 8411 44532 8430 44588
rect 8486 44532 8505 44588
rect 8411 44508 8505 44532
rect 8411 44452 8430 44508
rect 8486 44452 8505 44508
rect 8411 44428 8505 44452
rect 8411 44372 8430 44428
rect 8486 44372 8505 44428
rect 8411 44348 8505 44372
rect 8411 44292 8430 44348
rect 8486 44292 8505 44348
rect 8411 44264 8505 44292
rect 11301 44588 11395 44616
rect 11301 44532 11320 44588
rect 11376 44532 11395 44588
rect 11301 44508 11395 44532
rect 11301 44452 11320 44508
rect 11376 44452 11395 44508
rect 11301 44428 11395 44452
rect 11301 44372 11320 44428
rect 11376 44372 11395 44428
rect 11301 44348 11395 44372
rect 11301 44292 11320 44348
rect 11376 44292 11395 44348
rect 11301 44264 11395 44292
rect 14191 44588 14285 44616
rect 14191 44532 14210 44588
rect 14266 44532 14285 44588
rect 14191 44508 14285 44532
rect 14191 44452 14210 44508
rect 14266 44452 14285 44508
rect 14191 44428 14285 44452
rect 14191 44372 14210 44428
rect 14266 44372 14285 44428
rect 14191 44348 14285 44372
rect 14191 44292 14210 44348
rect 14266 44292 14285 44348
rect 14191 44264 14285 44292
rect 17081 44588 17175 44616
rect 17081 44532 17100 44588
rect 17156 44532 17175 44588
rect 17081 44508 17175 44532
rect 17081 44452 17100 44508
rect 17156 44452 17175 44508
rect 17081 44428 17175 44452
rect 17081 44372 17100 44428
rect 17156 44372 17175 44428
rect 17081 44348 17175 44372
rect 17081 44292 17100 44348
rect 17156 44292 17175 44348
rect 17081 44264 17175 44292
rect 19971 44588 20065 44616
rect 19971 44532 19990 44588
rect 20046 44532 20065 44588
rect 19971 44508 20065 44532
rect 19971 44452 19990 44508
rect 20046 44452 20065 44508
rect 19971 44428 20065 44452
rect 19971 44372 19990 44428
rect 20046 44372 20065 44428
rect 19971 44348 20065 44372
rect 19971 44292 19990 44348
rect 20046 44292 20065 44348
rect 19971 44264 20065 44292
rect 22861 44588 22955 44616
rect 22861 44532 22880 44588
rect 22936 44532 22955 44588
rect 22861 44508 22955 44532
rect 22861 44452 22880 44508
rect 22936 44452 22955 44508
rect 22861 44428 22955 44452
rect 22861 44372 22880 44428
rect 22936 44372 22955 44428
rect 22861 44348 22955 44372
rect 22861 44292 22880 44348
rect 22936 44292 22955 44348
rect 22861 44264 22955 44292
rect 25751 44588 25845 44616
rect 25751 44532 25770 44588
rect 25826 44532 25845 44588
rect 25751 44508 25845 44532
rect 25751 44452 25770 44508
rect 25826 44452 25845 44508
rect 25751 44428 25845 44452
rect 25751 44372 25770 44428
rect 25826 44372 25845 44428
rect 25751 44348 25845 44372
rect 25751 44292 25770 44348
rect 25826 44292 25845 44348
rect 25751 44264 25845 44292
rect 28641 44588 28735 44616
rect 28641 44532 28660 44588
rect 28716 44532 28735 44588
rect 28641 44508 28735 44532
rect 28641 44452 28660 44508
rect 28716 44452 28735 44508
rect 28641 44428 28735 44452
rect 28641 44372 28660 44428
rect 28716 44372 28735 44428
rect 28641 44348 28735 44372
rect 28641 44292 28660 44348
rect 28716 44292 28735 44348
rect 28641 44264 28735 44292
rect 31531 44588 31625 44616
rect 31531 44532 31550 44588
rect 31606 44532 31625 44588
rect 31531 44508 31625 44532
rect 31531 44452 31550 44508
rect 31606 44452 31625 44508
rect 31531 44428 31625 44452
rect 31531 44372 31550 44428
rect 31606 44372 31625 44428
rect 31531 44348 31625 44372
rect 31531 44292 31550 44348
rect 31606 44292 31625 44348
rect 31531 44264 31625 44292
rect 34421 44588 34515 44616
rect 34421 44532 34440 44588
rect 34496 44532 34515 44588
rect 34421 44508 34515 44532
rect 34421 44452 34440 44508
rect 34496 44452 34515 44508
rect 34421 44428 34515 44452
rect 34421 44372 34440 44428
rect 34496 44372 34515 44428
rect 34421 44348 34515 44372
rect 34421 44292 34440 44348
rect 34496 44292 34515 44348
rect 34421 44264 34515 44292
rect 37311 44588 37405 44616
rect 37311 44532 37330 44588
rect 37386 44532 37405 44588
rect 37311 44508 37405 44532
rect 37311 44452 37330 44508
rect 37386 44452 37405 44508
rect 37311 44428 37405 44452
rect 37311 44372 37330 44428
rect 37386 44372 37405 44428
rect 37311 44348 37405 44372
rect 37311 44292 37330 44348
rect 37386 44292 37405 44348
rect 37311 44264 37405 44292
rect 40201 44588 40295 44616
rect 40201 44532 40220 44588
rect 40276 44532 40295 44588
rect 40201 44508 40295 44532
rect 40201 44452 40220 44508
rect 40276 44452 40295 44508
rect 40201 44428 40295 44452
rect 40201 44372 40220 44428
rect 40276 44372 40295 44428
rect 40201 44348 40295 44372
rect 40201 44292 40220 44348
rect 40276 44292 40295 44348
rect 40201 44264 40295 44292
rect 43091 44588 43185 44616
rect 43091 44532 43110 44588
rect 43166 44532 43185 44588
rect 43091 44508 43185 44532
rect 43091 44452 43110 44508
rect 43166 44452 43185 44508
rect 43091 44428 43185 44452
rect 43091 44372 43110 44428
rect 43166 44372 43185 44428
rect 43091 44348 43185 44372
rect 43091 44292 43110 44348
rect 43166 44292 43185 44348
rect 43091 44264 43185 44292
rect 45981 44588 46075 44616
rect 45981 44532 46000 44588
rect 46056 44532 46075 44588
rect 45981 44508 46075 44532
rect 45981 44452 46000 44508
rect 46056 44452 46075 44508
rect 45981 44428 46075 44452
rect 45981 44372 46000 44428
rect 46056 44372 46075 44428
rect 45981 44348 46075 44372
rect 45981 44292 46000 44348
rect 46056 44292 46075 44348
rect 45981 44264 46075 44292
rect 52210 44588 52320 44616
rect 52210 44532 52237 44588
rect 52293 44532 52320 44588
rect 52210 44508 52320 44532
rect 52210 44452 52237 44508
rect 52293 44452 52320 44508
rect 52210 44428 52320 44452
rect 52210 44372 52237 44428
rect 52293 44372 52320 44428
rect 52210 44348 52320 44372
rect 52210 44292 52237 44348
rect 52293 44292 52320 44348
rect 52210 44264 52320 44292
rect 53602 44588 53730 44616
rect 53602 44532 53638 44588
rect 53694 44532 53730 44588
rect 53602 44508 53730 44532
rect 53602 44452 53638 44508
rect 53694 44452 53730 44508
rect 53602 44428 53730 44452
rect 53602 44372 53638 44428
rect 53694 44372 53730 44428
rect 53602 44348 53730 44372
rect 53602 44292 53638 44348
rect 53694 44292 53730 44348
rect 53602 44264 53730 44292
rect 54514 44588 54642 44616
rect 54514 44532 54550 44588
rect 54606 44532 54642 44588
rect 54514 44508 54642 44532
rect 54514 44452 54550 44508
rect 54606 44452 54642 44508
rect 54514 44428 54642 44452
rect 54514 44372 54550 44428
rect 54606 44372 54642 44428
rect 54514 44348 54642 44372
rect 54514 44292 54550 44348
rect 54606 44292 54642 44348
rect 54514 44264 54642 44292
rect 54910 44588 55026 44616
rect 54910 44532 54940 44588
rect 54996 44532 55026 44588
rect 54910 44508 55026 44532
rect 54910 44452 54940 44508
rect 54996 44452 55026 44508
rect 54910 44428 55026 44452
rect 54910 44372 54940 44428
rect 54996 44372 55026 44428
rect 54910 44348 55026 44372
rect 54910 44292 54940 44348
rect 54996 44292 55026 44348
rect 54910 44264 55026 44292
rect 55620 44588 55748 44616
rect 55620 44532 55656 44588
rect 55712 44532 55748 44588
rect 55620 44508 55748 44532
rect 55620 44452 55656 44508
rect 55712 44452 55748 44508
rect 55620 44428 55748 44452
rect 55620 44372 55656 44428
rect 55712 44372 55748 44428
rect 55620 44348 55748 44372
rect 55620 44292 55656 44348
rect 55712 44292 55748 44348
rect 55620 44264 55748 44292
rect 56198 44588 56326 44616
rect 56198 44532 56234 44588
rect 56290 44532 56326 44588
rect 56198 44508 56326 44532
rect 56198 44452 56234 44508
rect 56290 44452 56326 44508
rect 56198 44428 56326 44452
rect 56198 44372 56234 44428
rect 56290 44372 56326 44428
rect 56198 44348 56326 44372
rect 56198 44292 56234 44348
rect 56290 44292 56326 44348
rect 56198 44264 56326 44292
rect 56649 44588 56765 44616
rect 56649 44532 56679 44588
rect 56735 44532 56765 44588
rect 56649 44508 56765 44532
rect 56649 44452 56679 44508
rect 56735 44452 56765 44508
rect 56649 44428 56765 44452
rect 56649 44372 56679 44428
rect 56735 44372 56765 44428
rect 56649 44348 56765 44372
rect 56649 44292 56679 44348
rect 56735 44292 56765 44348
rect 56649 44264 56765 44292
rect 56953 44588 57069 44616
rect 56953 44532 56983 44588
rect 57039 44532 57069 44588
rect 56953 44508 57069 44532
rect 56953 44452 56983 44508
rect 57039 44452 57069 44508
rect 56953 44428 57069 44452
rect 56953 44372 56983 44428
rect 57039 44372 57069 44428
rect 56953 44348 57069 44372
rect 56953 44292 56983 44348
rect 57039 44292 57069 44348
rect 56953 44264 57069 44292
rect 57795 44588 57911 44616
rect 57795 44532 57825 44588
rect 57881 44532 57911 44588
rect 57795 44508 57911 44532
rect 57795 44452 57825 44508
rect 57881 44452 57911 44508
rect 57795 44428 57911 44452
rect 57795 44372 57825 44428
rect 57881 44372 57911 44428
rect 57795 44348 57911 44372
rect 57795 44292 57825 44348
rect 57881 44292 57911 44348
rect 57795 44264 57911 44292
rect 58345 44588 58409 44616
rect 58345 44532 58349 44588
rect 58405 44532 58409 44588
rect 58345 44508 58409 44532
rect 58345 44452 58349 44508
rect 58405 44452 58409 44508
rect 58345 44428 58409 44452
rect 58345 44372 58349 44428
rect 58405 44372 58409 44428
rect 58345 44348 58409 44372
rect 58345 44292 58349 44348
rect 58405 44292 58409 44348
rect 58345 44264 58409 44292
rect 59018 44588 59134 44616
rect 59018 44532 59048 44588
rect 59104 44532 59134 44588
rect 59018 44508 59134 44532
rect 59018 44452 59048 44508
rect 59104 44452 59134 44508
rect 59018 44428 59134 44452
rect 59018 44372 59048 44428
rect 59104 44372 59134 44428
rect 59018 44348 59134 44372
rect 59018 44292 59048 44348
rect 59104 44292 59134 44348
rect 59018 44264 59134 44292
rect 60296 44588 60412 44616
rect 60296 44532 60326 44588
rect 60382 44532 60412 44588
rect 60296 44508 60412 44532
rect 60296 44452 60326 44508
rect 60382 44452 60412 44508
rect 60296 44428 60412 44452
rect 60296 44372 60326 44428
rect 60382 44372 60412 44428
rect 60296 44348 60412 44372
rect 60296 44292 60326 44348
rect 60382 44292 60412 44348
rect 60296 44264 60412 44292
rect 60454 44588 60570 44616
rect 60454 44532 60484 44588
rect 60540 44532 60570 44588
rect 60454 44508 60570 44532
rect 60454 44452 60484 44508
rect 60540 44452 60570 44508
rect 60454 44428 60570 44452
rect 60454 44372 60484 44428
rect 60540 44372 60570 44428
rect 60454 44348 60570 44372
rect 60454 44292 60484 44348
rect 60540 44292 60570 44348
rect 60454 44264 60570 44292
rect 62509 44588 62683 44616
rect 62509 44532 62528 44588
rect 62584 44532 62608 44588
rect 62664 44532 62683 44588
rect 62509 44508 62683 44532
rect 62509 44452 62528 44508
rect 62584 44452 62608 44508
rect 62664 44452 62683 44508
rect 62509 44428 62683 44452
rect 62509 44372 62528 44428
rect 62584 44372 62608 44428
rect 62664 44372 62683 44428
rect 62509 44348 62683 44372
rect 62509 44292 62528 44348
rect 62584 44292 62608 44348
rect 62664 44292 62683 44348
rect 62509 44264 62683 44292
rect 2152 42236 2352 42264
rect 2152 42180 2184 42236
rect 2240 42180 2264 42236
rect 2320 42180 2352 42236
rect 2152 42156 2352 42180
rect 2152 42100 2184 42156
rect 2240 42100 2264 42156
rect 2320 42100 2352 42156
rect 2152 42076 2352 42100
rect 2152 42020 2184 42076
rect 2240 42020 2264 42076
rect 2320 42020 2352 42076
rect 2152 41996 2352 42020
rect 2152 41940 2184 41996
rect 2240 41940 2264 41996
rect 2320 41940 2352 41996
rect 2152 41912 2352 41940
rect 5374 42236 5468 42264
rect 5374 42180 5393 42236
rect 5449 42180 5468 42236
rect 5374 42156 5468 42180
rect 5374 42100 5393 42156
rect 5449 42100 5468 42156
rect 5374 42076 5468 42100
rect 5374 42020 5393 42076
rect 5449 42020 5468 42076
rect 5374 41996 5468 42020
rect 5374 41940 5393 41996
rect 5449 41940 5468 41996
rect 5374 41912 5468 41940
rect 8264 42236 8358 42264
rect 8264 42180 8283 42236
rect 8339 42180 8358 42236
rect 8264 42156 8358 42180
rect 8264 42100 8283 42156
rect 8339 42100 8358 42156
rect 8264 42076 8358 42100
rect 8264 42020 8283 42076
rect 8339 42020 8358 42076
rect 8264 41996 8358 42020
rect 8264 41940 8283 41996
rect 8339 41940 8358 41996
rect 8264 41912 8358 41940
rect 11154 42236 11248 42264
rect 11154 42180 11173 42236
rect 11229 42180 11248 42236
rect 11154 42156 11248 42180
rect 11154 42100 11173 42156
rect 11229 42100 11248 42156
rect 11154 42076 11248 42100
rect 11154 42020 11173 42076
rect 11229 42020 11248 42076
rect 11154 41996 11248 42020
rect 11154 41940 11173 41996
rect 11229 41940 11248 41996
rect 11154 41912 11248 41940
rect 14044 42236 14138 42264
rect 14044 42180 14063 42236
rect 14119 42180 14138 42236
rect 14044 42156 14138 42180
rect 14044 42100 14063 42156
rect 14119 42100 14138 42156
rect 14044 42076 14138 42100
rect 14044 42020 14063 42076
rect 14119 42020 14138 42076
rect 14044 41996 14138 42020
rect 14044 41940 14063 41996
rect 14119 41940 14138 41996
rect 14044 41912 14138 41940
rect 16934 42236 17028 42264
rect 16934 42180 16953 42236
rect 17009 42180 17028 42236
rect 16934 42156 17028 42180
rect 16934 42100 16953 42156
rect 17009 42100 17028 42156
rect 16934 42076 17028 42100
rect 16934 42020 16953 42076
rect 17009 42020 17028 42076
rect 16934 41996 17028 42020
rect 16934 41940 16953 41996
rect 17009 41940 17028 41996
rect 16934 41912 17028 41940
rect 19824 42236 19918 42264
rect 19824 42180 19843 42236
rect 19899 42180 19918 42236
rect 19824 42156 19918 42180
rect 19824 42100 19843 42156
rect 19899 42100 19918 42156
rect 19824 42076 19918 42100
rect 19824 42020 19843 42076
rect 19899 42020 19918 42076
rect 19824 41996 19918 42020
rect 19824 41940 19843 41996
rect 19899 41940 19918 41996
rect 19824 41912 19918 41940
rect 22714 42236 22808 42264
rect 22714 42180 22733 42236
rect 22789 42180 22808 42236
rect 22714 42156 22808 42180
rect 22714 42100 22733 42156
rect 22789 42100 22808 42156
rect 22714 42076 22808 42100
rect 22714 42020 22733 42076
rect 22789 42020 22808 42076
rect 22714 41996 22808 42020
rect 22714 41940 22733 41996
rect 22789 41940 22808 41996
rect 22714 41912 22808 41940
rect 25604 42236 25698 42264
rect 25604 42180 25623 42236
rect 25679 42180 25698 42236
rect 25604 42156 25698 42180
rect 25604 42100 25623 42156
rect 25679 42100 25698 42156
rect 25604 42076 25698 42100
rect 25604 42020 25623 42076
rect 25679 42020 25698 42076
rect 25604 41996 25698 42020
rect 25604 41940 25623 41996
rect 25679 41940 25698 41996
rect 25604 41912 25698 41940
rect 28494 42236 28588 42264
rect 28494 42180 28513 42236
rect 28569 42180 28588 42236
rect 28494 42156 28588 42180
rect 28494 42100 28513 42156
rect 28569 42100 28588 42156
rect 28494 42076 28588 42100
rect 28494 42020 28513 42076
rect 28569 42020 28588 42076
rect 28494 41996 28588 42020
rect 28494 41940 28513 41996
rect 28569 41940 28588 41996
rect 28494 41912 28588 41940
rect 31384 42236 31478 42264
rect 31384 42180 31403 42236
rect 31459 42180 31478 42236
rect 31384 42156 31478 42180
rect 31384 42100 31403 42156
rect 31459 42100 31478 42156
rect 31384 42076 31478 42100
rect 31384 42020 31403 42076
rect 31459 42020 31478 42076
rect 31384 41996 31478 42020
rect 31384 41940 31403 41996
rect 31459 41940 31478 41996
rect 31384 41912 31478 41940
rect 34274 42236 34368 42264
rect 34274 42180 34293 42236
rect 34349 42180 34368 42236
rect 34274 42156 34368 42180
rect 34274 42100 34293 42156
rect 34349 42100 34368 42156
rect 34274 42076 34368 42100
rect 34274 42020 34293 42076
rect 34349 42020 34368 42076
rect 34274 41996 34368 42020
rect 34274 41940 34293 41996
rect 34349 41940 34368 41996
rect 34274 41912 34368 41940
rect 37164 42236 37258 42264
rect 37164 42180 37183 42236
rect 37239 42180 37258 42236
rect 37164 42156 37258 42180
rect 37164 42100 37183 42156
rect 37239 42100 37258 42156
rect 37164 42076 37258 42100
rect 37164 42020 37183 42076
rect 37239 42020 37258 42076
rect 37164 41996 37258 42020
rect 37164 41940 37183 41996
rect 37239 41940 37258 41996
rect 37164 41912 37258 41940
rect 40054 42236 40148 42264
rect 40054 42180 40073 42236
rect 40129 42180 40148 42236
rect 40054 42156 40148 42180
rect 40054 42100 40073 42156
rect 40129 42100 40148 42156
rect 40054 42076 40148 42100
rect 40054 42020 40073 42076
rect 40129 42020 40148 42076
rect 40054 41996 40148 42020
rect 40054 41940 40073 41996
rect 40129 41940 40148 41996
rect 40054 41912 40148 41940
rect 42944 42236 43038 42264
rect 42944 42180 42963 42236
rect 43019 42180 43038 42236
rect 42944 42156 43038 42180
rect 42944 42100 42963 42156
rect 43019 42100 43038 42156
rect 42944 42076 43038 42100
rect 42944 42020 42963 42076
rect 43019 42020 43038 42076
rect 42944 41996 43038 42020
rect 42944 41940 42963 41996
rect 43019 41940 43038 41996
rect 42944 41912 43038 41940
rect 45834 42236 45928 42264
rect 45834 42180 45853 42236
rect 45909 42180 45928 42236
rect 45834 42156 45928 42180
rect 45834 42100 45853 42156
rect 45909 42100 45928 42156
rect 45834 42076 45928 42100
rect 45834 42020 45853 42076
rect 45909 42020 45928 42076
rect 45834 41996 45928 42020
rect 45834 41940 45853 41996
rect 45909 41940 45928 41996
rect 45834 41912 45928 41940
rect 48781 42236 48875 42264
rect 48781 42180 48800 42236
rect 48856 42180 48875 42236
rect 48781 42156 48875 42180
rect 48781 42100 48800 42156
rect 48856 42100 48875 42156
rect 48781 42076 48875 42100
rect 48781 42020 48800 42076
rect 48856 42020 48875 42076
rect 48781 41996 48875 42020
rect 48781 41940 48800 41996
rect 48856 41940 48875 41996
rect 48781 41912 48875 41940
rect 49630 42236 49830 42264
rect 49630 42180 49662 42236
rect 49718 42180 49742 42236
rect 49798 42180 49830 42236
rect 49630 42156 49830 42180
rect 49630 42100 49662 42156
rect 49718 42100 49742 42156
rect 49798 42100 49830 42156
rect 49630 42076 49830 42100
rect 49630 42020 49662 42076
rect 49718 42020 49742 42076
rect 49798 42020 49830 42076
rect 49630 41996 49830 42020
rect 49630 41940 49662 41996
rect 49718 41940 49742 41996
rect 49798 41940 49830 41996
rect 49630 41912 49830 41940
rect 52920 42236 53048 42264
rect 52920 42180 52956 42236
rect 53012 42180 53048 42236
rect 52920 42156 53048 42180
rect 52920 42100 52956 42156
rect 53012 42100 53048 42156
rect 52920 42076 53048 42100
rect 52920 42020 52956 42076
rect 53012 42020 53048 42076
rect 52920 41996 53048 42020
rect 52920 41940 52956 41996
rect 53012 41940 53048 41996
rect 52920 41912 53048 41940
rect 53078 42236 53206 42264
rect 53078 42180 53114 42236
rect 53170 42180 53206 42236
rect 53078 42156 53206 42180
rect 53078 42100 53114 42156
rect 53170 42100 53206 42156
rect 53078 42076 53206 42100
rect 53078 42020 53114 42076
rect 53170 42020 53206 42076
rect 53078 41996 53206 42020
rect 53078 41940 53114 41996
rect 53170 41940 53206 41996
rect 53078 41912 53206 41940
rect 53434 42236 53562 42264
rect 53434 42180 53470 42236
rect 53526 42180 53562 42236
rect 53434 42156 53562 42180
rect 53434 42100 53470 42156
rect 53526 42100 53562 42156
rect 53434 42076 53562 42100
rect 53434 42020 53470 42076
rect 53526 42020 53562 42076
rect 53434 41996 53562 42020
rect 53434 41940 53470 41996
rect 53526 41940 53562 41996
rect 53434 41912 53562 41940
rect 54752 42236 54880 42264
rect 54752 42180 54788 42236
rect 54844 42180 54880 42236
rect 54752 42156 54880 42180
rect 54752 42100 54788 42156
rect 54844 42100 54880 42156
rect 54752 42076 54880 42100
rect 54752 42020 54788 42076
rect 54844 42020 54880 42076
rect 54752 41996 54880 42020
rect 54752 41940 54788 41996
rect 54844 41940 54880 41996
rect 54752 41912 54880 41940
rect 55345 42236 55473 42264
rect 55345 42180 55381 42236
rect 55437 42180 55473 42236
rect 55345 42156 55473 42180
rect 55345 42100 55381 42156
rect 55437 42100 55473 42156
rect 55345 42076 55473 42100
rect 55345 42020 55381 42076
rect 55437 42020 55473 42076
rect 55345 41996 55473 42020
rect 55345 41940 55381 41996
rect 55437 41940 55473 41996
rect 55345 41912 55473 41940
rect 56491 42236 56619 42264
rect 56491 42180 56527 42236
rect 56583 42180 56619 42236
rect 56491 42156 56619 42180
rect 56491 42100 56527 42156
rect 56583 42100 56619 42156
rect 56491 42076 56619 42100
rect 56491 42020 56527 42076
rect 56583 42020 56619 42076
rect 56491 41996 56619 42020
rect 56491 41940 56527 41996
rect 56583 41940 56619 41996
rect 56491 41912 56619 41940
rect 57941 42236 58121 42264
rect 57941 42180 57963 42236
rect 58019 42180 58043 42236
rect 58099 42180 58121 42236
rect 57941 42156 58121 42180
rect 57941 42100 57963 42156
rect 58019 42100 58043 42156
rect 58099 42100 58121 42156
rect 57941 42076 58121 42100
rect 57941 42020 57963 42076
rect 58019 42020 58043 42076
rect 58099 42020 58121 42076
rect 57941 41996 58121 42020
rect 57941 41940 57963 41996
rect 58019 41940 58043 41996
rect 58099 41940 58121 41996
rect 57941 41912 58121 41940
rect 59164 42236 59304 42264
rect 59164 42180 59206 42236
rect 59262 42180 59304 42236
rect 59164 42156 59304 42180
rect 59164 42100 59206 42156
rect 59262 42100 59304 42156
rect 59164 42076 59304 42100
rect 59164 42020 59206 42076
rect 59262 42020 59304 42076
rect 59164 41996 59304 42020
rect 59164 41940 59206 41996
rect 59262 41940 59304 41996
rect 59164 41912 59304 41940
rect 59334 42236 59450 42264
rect 59334 42180 59364 42236
rect 59420 42180 59450 42236
rect 59334 42156 59450 42180
rect 59334 42100 59364 42156
rect 59420 42100 59450 42156
rect 59334 42076 59450 42100
rect 59334 42020 59364 42076
rect 59420 42020 59450 42076
rect 59334 41996 59450 42020
rect 59334 41940 59364 41996
rect 59420 41940 59450 41996
rect 59334 41912 59450 41940
rect 59642 42236 59758 42264
rect 59642 42180 59672 42236
rect 59728 42180 59758 42236
rect 59642 42156 59758 42180
rect 59642 42100 59672 42156
rect 59728 42100 59758 42156
rect 59642 42076 59758 42100
rect 59642 42020 59672 42076
rect 59728 42020 59758 42076
rect 59642 41996 59758 42020
rect 59642 41940 59672 41996
rect 59728 41940 59758 41996
rect 59642 41912 59758 41940
rect 59788 42236 59904 42264
rect 59788 42180 59818 42236
rect 59874 42180 59904 42236
rect 59788 42156 59904 42180
rect 59788 42100 59818 42156
rect 59874 42100 59904 42156
rect 59788 42076 59904 42100
rect 59788 42020 59818 42076
rect 59874 42020 59904 42076
rect 59788 41996 59904 42020
rect 59788 41940 59818 41996
rect 59874 41940 59904 41996
rect 59788 41912 59904 41940
rect 59934 42236 60110 42264
rect 59934 42180 59954 42236
rect 60010 42180 60034 42236
rect 60090 42180 60110 42236
rect 59934 42156 60110 42180
rect 59934 42100 59954 42156
rect 60010 42100 60034 42156
rect 60090 42100 60110 42156
rect 59934 42076 60110 42100
rect 59934 42020 59954 42076
rect 60010 42020 60034 42076
rect 60090 42020 60110 42076
rect 59934 41996 60110 42020
rect 59934 41940 59954 41996
rect 60010 41940 60034 41996
rect 60090 41940 60110 41996
rect 59934 41912 60110 41940
rect 62307 42236 62481 42264
rect 62307 42180 62326 42236
rect 62382 42180 62406 42236
rect 62462 42180 62481 42236
rect 62307 42156 62481 42180
rect 62307 42100 62326 42156
rect 62382 42100 62406 42156
rect 62462 42100 62481 42156
rect 62307 42076 62481 42100
rect 62307 42020 62326 42076
rect 62382 42020 62406 42076
rect 62462 42020 62481 42076
rect 62307 41996 62481 42020
rect 62307 41940 62326 41996
rect 62382 41940 62406 41996
rect 62462 41940 62481 41996
rect 62307 41912 62481 41940
rect 2020 34588 2124 34616
rect 2020 34532 2044 34588
rect 2100 34532 2124 34588
rect 2020 34508 2124 34532
rect 2020 34452 2044 34508
rect 2100 34452 2124 34508
rect 2020 34428 2124 34452
rect 2020 34372 2044 34428
rect 2100 34372 2124 34428
rect 2020 34348 2124 34372
rect 2020 34292 2044 34348
rect 2100 34292 2124 34348
rect 2020 34264 2124 34292
rect 5521 34588 5615 34616
rect 5521 34532 5540 34588
rect 5596 34532 5615 34588
rect 5521 34508 5615 34532
rect 5521 34452 5540 34508
rect 5596 34452 5615 34508
rect 5521 34428 5615 34452
rect 5521 34372 5540 34428
rect 5596 34372 5615 34428
rect 5521 34348 5615 34372
rect 5521 34292 5540 34348
rect 5596 34292 5615 34348
rect 5521 34264 5615 34292
rect 8411 34588 8505 34616
rect 8411 34532 8430 34588
rect 8486 34532 8505 34588
rect 8411 34508 8505 34532
rect 8411 34452 8430 34508
rect 8486 34452 8505 34508
rect 8411 34428 8505 34452
rect 8411 34372 8430 34428
rect 8486 34372 8505 34428
rect 8411 34348 8505 34372
rect 8411 34292 8430 34348
rect 8486 34292 8505 34348
rect 8411 34264 8505 34292
rect 11301 34588 11395 34616
rect 11301 34532 11320 34588
rect 11376 34532 11395 34588
rect 11301 34508 11395 34532
rect 11301 34452 11320 34508
rect 11376 34452 11395 34508
rect 11301 34428 11395 34452
rect 11301 34372 11320 34428
rect 11376 34372 11395 34428
rect 11301 34348 11395 34372
rect 11301 34292 11320 34348
rect 11376 34292 11395 34348
rect 11301 34264 11395 34292
rect 14191 34588 14285 34616
rect 14191 34532 14210 34588
rect 14266 34532 14285 34588
rect 14191 34508 14285 34532
rect 14191 34452 14210 34508
rect 14266 34452 14285 34508
rect 14191 34428 14285 34452
rect 14191 34372 14210 34428
rect 14266 34372 14285 34428
rect 14191 34348 14285 34372
rect 14191 34292 14210 34348
rect 14266 34292 14285 34348
rect 14191 34264 14285 34292
rect 17081 34588 17175 34616
rect 17081 34532 17100 34588
rect 17156 34532 17175 34588
rect 17081 34508 17175 34532
rect 17081 34452 17100 34508
rect 17156 34452 17175 34508
rect 17081 34428 17175 34452
rect 17081 34372 17100 34428
rect 17156 34372 17175 34428
rect 17081 34348 17175 34372
rect 17081 34292 17100 34348
rect 17156 34292 17175 34348
rect 17081 34264 17175 34292
rect 19971 34588 20065 34616
rect 19971 34532 19990 34588
rect 20046 34532 20065 34588
rect 19971 34508 20065 34532
rect 19971 34452 19990 34508
rect 20046 34452 20065 34508
rect 19971 34428 20065 34452
rect 19971 34372 19990 34428
rect 20046 34372 20065 34428
rect 19971 34348 20065 34372
rect 19971 34292 19990 34348
rect 20046 34292 20065 34348
rect 19971 34264 20065 34292
rect 22861 34588 22955 34616
rect 22861 34532 22880 34588
rect 22936 34532 22955 34588
rect 22861 34508 22955 34532
rect 22861 34452 22880 34508
rect 22936 34452 22955 34508
rect 22861 34428 22955 34452
rect 22861 34372 22880 34428
rect 22936 34372 22955 34428
rect 22861 34348 22955 34372
rect 22861 34292 22880 34348
rect 22936 34292 22955 34348
rect 22861 34264 22955 34292
rect 25751 34588 25845 34616
rect 25751 34532 25770 34588
rect 25826 34532 25845 34588
rect 25751 34508 25845 34532
rect 25751 34452 25770 34508
rect 25826 34452 25845 34508
rect 25751 34428 25845 34452
rect 25751 34372 25770 34428
rect 25826 34372 25845 34428
rect 25751 34348 25845 34372
rect 25751 34292 25770 34348
rect 25826 34292 25845 34348
rect 25751 34264 25845 34292
rect 28641 34588 28735 34616
rect 28641 34532 28660 34588
rect 28716 34532 28735 34588
rect 28641 34508 28735 34532
rect 28641 34452 28660 34508
rect 28716 34452 28735 34508
rect 28641 34428 28735 34452
rect 28641 34372 28660 34428
rect 28716 34372 28735 34428
rect 28641 34348 28735 34372
rect 28641 34292 28660 34348
rect 28716 34292 28735 34348
rect 28641 34264 28735 34292
rect 31531 34588 31625 34616
rect 31531 34532 31550 34588
rect 31606 34532 31625 34588
rect 31531 34508 31625 34532
rect 31531 34452 31550 34508
rect 31606 34452 31625 34508
rect 31531 34428 31625 34452
rect 31531 34372 31550 34428
rect 31606 34372 31625 34428
rect 31531 34348 31625 34372
rect 31531 34292 31550 34348
rect 31606 34292 31625 34348
rect 31531 34264 31625 34292
rect 34421 34588 34515 34616
rect 34421 34532 34440 34588
rect 34496 34532 34515 34588
rect 34421 34508 34515 34532
rect 34421 34452 34440 34508
rect 34496 34452 34515 34508
rect 34421 34428 34515 34452
rect 34421 34372 34440 34428
rect 34496 34372 34515 34428
rect 34421 34348 34515 34372
rect 34421 34292 34440 34348
rect 34496 34292 34515 34348
rect 34421 34264 34515 34292
rect 37311 34588 37405 34616
rect 37311 34532 37330 34588
rect 37386 34532 37405 34588
rect 37311 34508 37405 34532
rect 37311 34452 37330 34508
rect 37386 34452 37405 34508
rect 37311 34428 37405 34452
rect 37311 34372 37330 34428
rect 37386 34372 37405 34428
rect 37311 34348 37405 34372
rect 37311 34292 37330 34348
rect 37386 34292 37405 34348
rect 37311 34264 37405 34292
rect 40201 34588 40295 34616
rect 40201 34532 40220 34588
rect 40276 34532 40295 34588
rect 40201 34508 40295 34532
rect 40201 34452 40220 34508
rect 40276 34452 40295 34508
rect 40201 34428 40295 34452
rect 40201 34372 40220 34428
rect 40276 34372 40295 34428
rect 40201 34348 40295 34372
rect 40201 34292 40220 34348
rect 40276 34292 40295 34348
rect 40201 34264 40295 34292
rect 43091 34588 43185 34616
rect 43091 34532 43110 34588
rect 43166 34532 43185 34588
rect 43091 34508 43185 34532
rect 43091 34452 43110 34508
rect 43166 34452 43185 34508
rect 43091 34428 43185 34452
rect 43091 34372 43110 34428
rect 43166 34372 43185 34428
rect 43091 34348 43185 34372
rect 43091 34292 43110 34348
rect 43166 34292 43185 34348
rect 43091 34264 43185 34292
rect 45981 34588 46075 34616
rect 45981 34532 46000 34588
rect 46056 34532 46075 34588
rect 45981 34508 46075 34532
rect 45981 34452 46000 34508
rect 46056 34452 46075 34508
rect 45981 34428 46075 34452
rect 45981 34372 46000 34428
rect 46056 34372 46075 34428
rect 45981 34348 46075 34372
rect 45981 34292 46000 34348
rect 46056 34292 46075 34348
rect 45981 34264 46075 34292
rect 48989 34588 49083 34616
rect 48989 34532 49008 34588
rect 49064 34532 49083 34588
rect 48989 34508 49083 34532
rect 48989 34452 49008 34508
rect 49064 34452 49083 34508
rect 48989 34428 49083 34452
rect 48989 34372 49008 34428
rect 49064 34372 49083 34428
rect 48989 34348 49083 34372
rect 48989 34292 49008 34348
rect 49064 34292 49083 34348
rect 48989 34264 49083 34292
rect 52210 34588 52320 34616
rect 52210 34532 52237 34588
rect 52293 34532 52320 34588
rect 52210 34508 52320 34532
rect 52210 34452 52237 34508
rect 52293 34452 52320 34508
rect 52210 34428 52320 34452
rect 52210 34372 52237 34428
rect 52293 34372 52320 34428
rect 52210 34348 52320 34372
rect 52210 34292 52237 34348
rect 52293 34292 52320 34348
rect 52210 34264 52320 34292
rect 53602 34588 53730 34616
rect 53602 34532 53638 34588
rect 53694 34532 53730 34588
rect 53602 34508 53730 34532
rect 53602 34452 53638 34508
rect 53694 34452 53730 34508
rect 53602 34428 53730 34452
rect 53602 34372 53638 34428
rect 53694 34372 53730 34428
rect 53602 34348 53730 34372
rect 53602 34292 53638 34348
rect 53694 34292 53730 34348
rect 53602 34264 53730 34292
rect 53770 34588 53898 34616
rect 53770 34532 53806 34588
rect 53862 34532 53898 34588
rect 53770 34508 53898 34532
rect 53770 34452 53806 34508
rect 53862 34452 53898 34508
rect 53770 34428 53898 34452
rect 53770 34372 53806 34428
rect 53862 34372 53898 34428
rect 53770 34348 53898 34372
rect 53770 34292 53806 34348
rect 53862 34292 53898 34348
rect 53770 34264 53898 34292
rect 54514 34588 54642 34616
rect 54514 34532 54550 34588
rect 54606 34532 54642 34588
rect 54514 34508 54642 34532
rect 54514 34452 54550 34508
rect 54606 34452 54642 34508
rect 54514 34428 54642 34452
rect 54514 34372 54550 34428
rect 54606 34372 54642 34428
rect 54514 34348 54642 34372
rect 54514 34292 54550 34348
rect 54606 34292 54642 34348
rect 54514 34264 54642 34292
rect 54910 34588 55026 34616
rect 54910 34532 54940 34588
rect 54996 34532 55026 34588
rect 54910 34508 55026 34532
rect 54910 34452 54940 34508
rect 54996 34452 55026 34508
rect 54910 34428 55026 34452
rect 54910 34372 54940 34428
rect 54996 34372 55026 34428
rect 54910 34348 55026 34372
rect 54910 34292 54940 34348
rect 54996 34292 55026 34348
rect 54910 34264 55026 34292
rect 55620 34588 55748 34616
rect 55620 34532 55656 34588
rect 55712 34532 55748 34588
rect 55620 34508 55748 34532
rect 55620 34452 55656 34508
rect 55712 34452 55748 34508
rect 55620 34428 55748 34452
rect 55620 34372 55656 34428
rect 55712 34372 55748 34428
rect 55620 34348 55748 34372
rect 55620 34292 55656 34348
rect 55712 34292 55748 34348
rect 55620 34264 55748 34292
rect 56198 34588 56326 34616
rect 56198 34532 56234 34588
rect 56290 34532 56326 34588
rect 56198 34508 56326 34532
rect 56198 34452 56234 34508
rect 56290 34452 56326 34508
rect 56198 34428 56326 34452
rect 56198 34372 56234 34428
rect 56290 34372 56326 34428
rect 56198 34348 56326 34372
rect 56198 34292 56234 34348
rect 56290 34292 56326 34348
rect 56198 34264 56326 34292
rect 56649 34588 56765 34616
rect 56649 34532 56679 34588
rect 56735 34532 56765 34588
rect 56649 34508 56765 34532
rect 56649 34452 56679 34508
rect 56735 34452 56765 34508
rect 56649 34428 56765 34452
rect 56649 34372 56679 34428
rect 56735 34372 56765 34428
rect 56649 34348 56765 34372
rect 56649 34292 56679 34348
rect 56735 34292 56765 34348
rect 56649 34264 56765 34292
rect 56953 34588 57069 34616
rect 56953 34532 56983 34588
rect 57039 34532 57069 34588
rect 56953 34508 57069 34532
rect 56953 34452 56983 34508
rect 57039 34452 57069 34508
rect 56953 34428 57069 34452
rect 56953 34372 56983 34428
rect 57039 34372 57069 34428
rect 56953 34348 57069 34372
rect 56953 34292 56983 34348
rect 57039 34292 57069 34348
rect 56953 34264 57069 34292
rect 57795 34588 57911 34616
rect 57795 34532 57825 34588
rect 57881 34532 57911 34588
rect 57795 34508 57911 34532
rect 57795 34452 57825 34508
rect 57881 34452 57911 34508
rect 57795 34428 57911 34452
rect 57795 34372 57825 34428
rect 57881 34372 57911 34428
rect 57795 34348 57911 34372
rect 57795 34292 57825 34348
rect 57881 34292 57911 34348
rect 57795 34264 57911 34292
rect 58461 34588 58525 34616
rect 58461 34532 58465 34588
rect 58521 34532 58525 34588
rect 58461 34508 58525 34532
rect 58461 34452 58465 34508
rect 58521 34452 58525 34508
rect 58461 34428 58525 34452
rect 58461 34372 58465 34428
rect 58521 34372 58525 34428
rect 58461 34348 58525 34372
rect 58461 34292 58465 34348
rect 58521 34292 58525 34348
rect 58461 34264 58525 34292
rect 59018 34588 59134 34616
rect 59018 34532 59048 34588
rect 59104 34532 59134 34588
rect 59018 34508 59134 34532
rect 59018 34452 59048 34508
rect 59104 34452 59134 34508
rect 59018 34428 59134 34452
rect 59018 34372 59048 34428
rect 59104 34372 59134 34428
rect 59018 34348 59134 34372
rect 59018 34292 59048 34348
rect 59104 34292 59134 34348
rect 59018 34264 59134 34292
rect 60296 34588 60412 34616
rect 60296 34532 60326 34588
rect 60382 34532 60412 34588
rect 60296 34508 60412 34532
rect 60296 34452 60326 34508
rect 60382 34452 60412 34508
rect 60296 34428 60412 34452
rect 60296 34372 60326 34428
rect 60382 34372 60412 34428
rect 60296 34348 60412 34372
rect 60296 34292 60326 34348
rect 60382 34292 60412 34348
rect 60296 34264 60412 34292
rect 60454 34588 60570 34616
rect 60454 34532 60484 34588
rect 60540 34532 60570 34588
rect 60454 34508 60570 34532
rect 60454 34452 60484 34508
rect 60540 34452 60570 34508
rect 60454 34428 60570 34452
rect 60454 34372 60484 34428
rect 60540 34372 60570 34428
rect 60454 34348 60570 34372
rect 60454 34292 60484 34348
rect 60540 34292 60570 34348
rect 60454 34264 60570 34292
rect 62509 34588 62683 34616
rect 62509 34532 62528 34588
rect 62584 34532 62608 34588
rect 62664 34532 62683 34588
rect 62509 34508 62683 34532
rect 62509 34452 62528 34508
rect 62584 34452 62608 34508
rect 62664 34452 62683 34508
rect 62509 34428 62683 34452
rect 62509 34372 62528 34428
rect 62584 34372 62608 34428
rect 62664 34372 62683 34428
rect 62509 34348 62683 34372
rect 62509 34292 62528 34348
rect 62584 34292 62608 34348
rect 62664 34292 62683 34348
rect 62509 34264 62683 34292
rect 2152 32236 2352 32264
rect 2152 32180 2184 32236
rect 2240 32180 2264 32236
rect 2320 32180 2352 32236
rect 2152 32156 2352 32180
rect 2152 32100 2184 32156
rect 2240 32100 2264 32156
rect 2320 32100 2352 32156
rect 2152 32076 2352 32100
rect 2152 32020 2184 32076
rect 2240 32020 2264 32076
rect 2320 32020 2352 32076
rect 2152 31996 2352 32020
rect 2152 31940 2184 31996
rect 2240 31940 2264 31996
rect 2320 31940 2352 31996
rect 2152 31912 2352 31940
rect 5374 32236 5468 32264
rect 5374 32180 5393 32236
rect 5449 32180 5468 32236
rect 5374 32156 5468 32180
rect 5374 32100 5393 32156
rect 5449 32100 5468 32156
rect 5374 32076 5468 32100
rect 5374 32020 5393 32076
rect 5449 32020 5468 32076
rect 5374 31996 5468 32020
rect 5374 31940 5393 31996
rect 5449 31940 5468 31996
rect 5374 31912 5468 31940
rect 8264 32236 8358 32264
rect 8264 32180 8283 32236
rect 8339 32180 8358 32236
rect 8264 32156 8358 32180
rect 8264 32100 8283 32156
rect 8339 32100 8358 32156
rect 8264 32076 8358 32100
rect 8264 32020 8283 32076
rect 8339 32020 8358 32076
rect 8264 31996 8358 32020
rect 8264 31940 8283 31996
rect 8339 31940 8358 31996
rect 8264 31912 8358 31940
rect 11154 32236 11248 32264
rect 11154 32180 11173 32236
rect 11229 32180 11248 32236
rect 11154 32156 11248 32180
rect 11154 32100 11173 32156
rect 11229 32100 11248 32156
rect 11154 32076 11248 32100
rect 11154 32020 11173 32076
rect 11229 32020 11248 32076
rect 11154 31996 11248 32020
rect 11154 31940 11173 31996
rect 11229 31940 11248 31996
rect 11154 31912 11248 31940
rect 14044 32236 14138 32264
rect 14044 32180 14063 32236
rect 14119 32180 14138 32236
rect 14044 32156 14138 32180
rect 14044 32100 14063 32156
rect 14119 32100 14138 32156
rect 14044 32076 14138 32100
rect 14044 32020 14063 32076
rect 14119 32020 14138 32076
rect 14044 31996 14138 32020
rect 14044 31940 14063 31996
rect 14119 31940 14138 31996
rect 14044 31912 14138 31940
rect 16934 32236 17028 32264
rect 16934 32180 16953 32236
rect 17009 32180 17028 32236
rect 16934 32156 17028 32180
rect 16934 32100 16953 32156
rect 17009 32100 17028 32156
rect 16934 32076 17028 32100
rect 16934 32020 16953 32076
rect 17009 32020 17028 32076
rect 16934 31996 17028 32020
rect 16934 31940 16953 31996
rect 17009 31940 17028 31996
rect 16934 31912 17028 31940
rect 19824 32236 19918 32264
rect 19824 32180 19843 32236
rect 19899 32180 19918 32236
rect 19824 32156 19918 32180
rect 19824 32100 19843 32156
rect 19899 32100 19918 32156
rect 19824 32076 19918 32100
rect 19824 32020 19843 32076
rect 19899 32020 19918 32076
rect 19824 31996 19918 32020
rect 19824 31940 19843 31996
rect 19899 31940 19918 31996
rect 19824 31912 19918 31940
rect 22714 32236 22808 32264
rect 22714 32180 22733 32236
rect 22789 32180 22808 32236
rect 22714 32156 22808 32180
rect 22714 32100 22733 32156
rect 22789 32100 22808 32156
rect 22714 32076 22808 32100
rect 22714 32020 22733 32076
rect 22789 32020 22808 32076
rect 22714 31996 22808 32020
rect 22714 31940 22733 31996
rect 22789 31940 22808 31996
rect 22714 31912 22808 31940
rect 25604 32236 25698 32264
rect 25604 32180 25623 32236
rect 25679 32180 25698 32236
rect 25604 32156 25698 32180
rect 25604 32100 25623 32156
rect 25679 32100 25698 32156
rect 25604 32076 25698 32100
rect 25604 32020 25623 32076
rect 25679 32020 25698 32076
rect 25604 31996 25698 32020
rect 25604 31940 25623 31996
rect 25679 31940 25698 31996
rect 25604 31912 25698 31940
rect 28494 32236 28588 32264
rect 28494 32180 28513 32236
rect 28569 32180 28588 32236
rect 28494 32156 28588 32180
rect 28494 32100 28513 32156
rect 28569 32100 28588 32156
rect 28494 32076 28588 32100
rect 28494 32020 28513 32076
rect 28569 32020 28588 32076
rect 28494 31996 28588 32020
rect 28494 31940 28513 31996
rect 28569 31940 28588 31996
rect 28494 31912 28588 31940
rect 31384 32236 31478 32264
rect 31384 32180 31403 32236
rect 31459 32180 31478 32236
rect 31384 32156 31478 32180
rect 31384 32100 31403 32156
rect 31459 32100 31478 32156
rect 31384 32076 31478 32100
rect 31384 32020 31403 32076
rect 31459 32020 31478 32076
rect 31384 31996 31478 32020
rect 31384 31940 31403 31996
rect 31459 31940 31478 31996
rect 31384 31912 31478 31940
rect 34274 32236 34368 32264
rect 34274 32180 34293 32236
rect 34349 32180 34368 32236
rect 34274 32156 34368 32180
rect 34274 32100 34293 32156
rect 34349 32100 34368 32156
rect 34274 32076 34368 32100
rect 34274 32020 34293 32076
rect 34349 32020 34368 32076
rect 34274 31996 34368 32020
rect 34274 31940 34293 31996
rect 34349 31940 34368 31996
rect 34274 31912 34368 31940
rect 37164 32236 37258 32264
rect 37164 32180 37183 32236
rect 37239 32180 37258 32236
rect 37164 32156 37258 32180
rect 37164 32100 37183 32156
rect 37239 32100 37258 32156
rect 37164 32076 37258 32100
rect 37164 32020 37183 32076
rect 37239 32020 37258 32076
rect 37164 31996 37258 32020
rect 37164 31940 37183 31996
rect 37239 31940 37258 31996
rect 37164 31912 37258 31940
rect 40054 32236 40148 32264
rect 40054 32180 40073 32236
rect 40129 32180 40148 32236
rect 40054 32156 40148 32180
rect 40054 32100 40073 32156
rect 40129 32100 40148 32156
rect 40054 32076 40148 32100
rect 40054 32020 40073 32076
rect 40129 32020 40148 32076
rect 40054 31996 40148 32020
rect 40054 31940 40073 31996
rect 40129 31940 40148 31996
rect 40054 31912 40148 31940
rect 42944 32236 43038 32264
rect 42944 32180 42963 32236
rect 43019 32180 43038 32236
rect 42944 32156 43038 32180
rect 42944 32100 42963 32156
rect 43019 32100 43038 32156
rect 42944 32076 43038 32100
rect 42944 32020 42963 32076
rect 43019 32020 43038 32076
rect 42944 31996 43038 32020
rect 42944 31940 42963 31996
rect 43019 31940 43038 31996
rect 42944 31912 43038 31940
rect 45834 32236 45928 32264
rect 45834 32180 45853 32236
rect 45909 32180 45928 32236
rect 45834 32156 45928 32180
rect 45834 32100 45853 32156
rect 45909 32100 45928 32156
rect 45834 32076 45928 32100
rect 45834 32020 45853 32076
rect 45909 32020 45928 32076
rect 45834 31996 45928 32020
rect 45834 31940 45853 31996
rect 45909 31940 45928 31996
rect 45834 31912 45928 31940
rect 48781 32236 48875 32264
rect 48781 32180 48800 32236
rect 48856 32180 48875 32236
rect 48781 32156 48875 32180
rect 48781 32100 48800 32156
rect 48856 32100 48875 32156
rect 48781 32076 48875 32100
rect 48781 32020 48800 32076
rect 48856 32020 48875 32076
rect 48781 31996 48875 32020
rect 48781 31940 48800 31996
rect 48856 31940 48875 31996
rect 48781 31912 48875 31940
rect 49630 32236 49830 32264
rect 49630 32180 49662 32236
rect 49718 32180 49742 32236
rect 49798 32180 49830 32236
rect 49630 32156 49830 32180
rect 49630 32100 49662 32156
rect 49718 32100 49742 32156
rect 49798 32100 49830 32156
rect 49630 32076 49830 32100
rect 49630 32020 49662 32076
rect 49718 32020 49742 32076
rect 49798 32020 49830 32076
rect 49630 31996 49830 32020
rect 49630 31940 49662 31996
rect 49718 31940 49742 31996
rect 49798 31940 49830 31996
rect 49630 31912 49830 31940
rect 52920 32236 53048 32264
rect 52920 32180 52956 32236
rect 53012 32180 53048 32236
rect 52920 32156 53048 32180
rect 52920 32100 52956 32156
rect 53012 32100 53048 32156
rect 52920 32076 53048 32100
rect 52920 32020 52956 32076
rect 53012 32020 53048 32076
rect 52920 31996 53048 32020
rect 52920 31940 52956 31996
rect 53012 31940 53048 31996
rect 52920 31912 53048 31940
rect 53078 32236 53206 32264
rect 53078 32180 53114 32236
rect 53170 32180 53206 32236
rect 53078 32156 53206 32180
rect 53078 32100 53114 32156
rect 53170 32100 53206 32156
rect 53078 32076 53206 32100
rect 53078 32020 53114 32076
rect 53170 32020 53206 32076
rect 53078 31996 53206 32020
rect 53078 31940 53114 31996
rect 53170 31940 53206 31996
rect 53078 31912 53206 31940
rect 53434 32236 53562 32264
rect 53434 32180 53470 32236
rect 53526 32180 53562 32236
rect 53434 32156 53562 32180
rect 53434 32100 53470 32156
rect 53526 32100 53562 32156
rect 53434 32076 53562 32100
rect 53434 32020 53470 32076
rect 53526 32020 53562 32076
rect 53434 31996 53562 32020
rect 53434 31940 53470 31996
rect 53526 31940 53562 31996
rect 53434 31912 53562 31940
rect 54752 32236 54880 32264
rect 54752 32180 54788 32236
rect 54844 32180 54880 32236
rect 54752 32156 54880 32180
rect 54752 32100 54788 32156
rect 54844 32100 54880 32156
rect 54752 32076 54880 32100
rect 54752 32020 54788 32076
rect 54844 32020 54880 32076
rect 54752 31996 54880 32020
rect 54752 31940 54788 31996
rect 54844 31940 54880 31996
rect 54752 31912 54880 31940
rect 55345 32236 55473 32264
rect 55345 32180 55381 32236
rect 55437 32180 55473 32236
rect 55345 32156 55473 32180
rect 55345 32100 55381 32156
rect 55437 32100 55473 32156
rect 55345 32076 55473 32100
rect 55345 32020 55381 32076
rect 55437 32020 55473 32076
rect 55345 31996 55473 32020
rect 55345 31940 55381 31996
rect 55437 31940 55473 31996
rect 55345 31912 55473 31940
rect 56491 32236 56619 32264
rect 56491 32180 56527 32236
rect 56583 32180 56619 32236
rect 56491 32156 56619 32180
rect 56491 32100 56527 32156
rect 56583 32100 56619 32156
rect 56491 32076 56619 32100
rect 56491 32020 56527 32076
rect 56583 32020 56619 32076
rect 56491 31996 56619 32020
rect 56491 31940 56527 31996
rect 56583 31940 56619 31996
rect 56491 31912 56619 31940
rect 57941 32236 58121 32264
rect 57941 32180 57963 32236
rect 58019 32180 58043 32236
rect 58099 32180 58121 32236
rect 57941 32156 58121 32180
rect 57941 32100 57963 32156
rect 58019 32100 58043 32156
rect 58099 32100 58121 32156
rect 57941 32076 58121 32100
rect 57941 32020 57963 32076
rect 58019 32020 58043 32076
rect 58099 32020 58121 32076
rect 57941 31996 58121 32020
rect 57941 31940 57963 31996
rect 58019 31940 58043 31996
rect 58099 31940 58121 31996
rect 57941 31912 58121 31940
rect 59164 32236 59304 32264
rect 59164 32180 59206 32236
rect 59262 32180 59304 32236
rect 59164 32156 59304 32180
rect 59164 32100 59206 32156
rect 59262 32100 59304 32156
rect 59164 32076 59304 32100
rect 59164 32020 59206 32076
rect 59262 32020 59304 32076
rect 59164 31996 59304 32020
rect 59164 31940 59206 31996
rect 59262 31940 59304 31996
rect 59164 31912 59304 31940
rect 59334 32236 59450 32264
rect 59334 32180 59364 32236
rect 59420 32180 59450 32236
rect 59334 32156 59450 32180
rect 59334 32100 59364 32156
rect 59420 32100 59450 32156
rect 59334 32076 59450 32100
rect 59334 32020 59364 32076
rect 59420 32020 59450 32076
rect 59334 31996 59450 32020
rect 59334 31940 59364 31996
rect 59420 31940 59450 31996
rect 59334 31912 59450 31940
rect 59642 32236 59758 32264
rect 59642 32180 59672 32236
rect 59728 32180 59758 32236
rect 59642 32156 59758 32180
rect 59642 32100 59672 32156
rect 59728 32100 59758 32156
rect 59642 32076 59758 32100
rect 59642 32020 59672 32076
rect 59728 32020 59758 32076
rect 59642 31996 59758 32020
rect 59642 31940 59672 31996
rect 59728 31940 59758 31996
rect 59642 31912 59758 31940
rect 59788 32236 59904 32264
rect 59788 32180 59818 32236
rect 59874 32180 59904 32236
rect 59788 32156 59904 32180
rect 59788 32100 59818 32156
rect 59874 32100 59904 32156
rect 59788 32076 59904 32100
rect 59788 32020 59818 32076
rect 59874 32020 59904 32076
rect 59788 31996 59904 32020
rect 59788 31940 59818 31996
rect 59874 31940 59904 31996
rect 59788 31912 59904 31940
rect 59934 32236 60110 32264
rect 59934 32180 59954 32236
rect 60010 32180 60034 32236
rect 60090 32180 60110 32236
rect 59934 32156 60110 32180
rect 59934 32100 59954 32156
rect 60010 32100 60034 32156
rect 60090 32100 60110 32156
rect 59934 32076 60110 32100
rect 59934 32020 59954 32076
rect 60010 32020 60034 32076
rect 60090 32020 60110 32076
rect 59934 31996 60110 32020
rect 59934 31940 59954 31996
rect 60010 31940 60034 31996
rect 60090 31940 60110 31996
rect 59934 31912 60110 31940
rect 62307 32236 62481 32264
rect 62307 32180 62326 32236
rect 62382 32180 62406 32236
rect 62462 32180 62481 32236
rect 62307 32156 62481 32180
rect 62307 32100 62326 32156
rect 62382 32100 62406 32156
rect 62462 32100 62481 32156
rect 62307 32076 62481 32100
rect 62307 32020 62326 32076
rect 62382 32020 62406 32076
rect 62462 32020 62481 32076
rect 62307 31996 62481 32020
rect 62307 31940 62326 31996
rect 62382 31940 62406 31996
rect 62462 31940 62481 31996
rect 62307 31912 62481 31940
rect 2020 24588 2124 24616
rect 2020 24532 2044 24588
rect 2100 24532 2124 24588
rect 2020 24508 2124 24532
rect 2020 24452 2044 24508
rect 2100 24452 2124 24508
rect 2020 24428 2124 24452
rect 2020 24372 2044 24428
rect 2100 24372 2124 24428
rect 2020 24348 2124 24372
rect 2020 24292 2044 24348
rect 2100 24292 2124 24348
rect 2020 24264 2124 24292
rect 5521 24588 5615 24616
rect 5521 24532 5540 24588
rect 5596 24532 5615 24588
rect 5521 24508 5615 24532
rect 5521 24452 5540 24508
rect 5596 24452 5615 24508
rect 5521 24428 5615 24452
rect 5521 24372 5540 24428
rect 5596 24372 5615 24428
rect 5521 24348 5615 24372
rect 5521 24292 5540 24348
rect 5596 24292 5615 24348
rect 5521 24264 5615 24292
rect 8411 24588 8505 24616
rect 8411 24532 8430 24588
rect 8486 24532 8505 24588
rect 8411 24508 8505 24532
rect 8411 24452 8430 24508
rect 8486 24452 8505 24508
rect 8411 24428 8505 24452
rect 8411 24372 8430 24428
rect 8486 24372 8505 24428
rect 8411 24348 8505 24372
rect 8411 24292 8430 24348
rect 8486 24292 8505 24348
rect 8411 24264 8505 24292
rect 11301 24588 11395 24616
rect 11301 24532 11320 24588
rect 11376 24532 11395 24588
rect 11301 24508 11395 24532
rect 11301 24452 11320 24508
rect 11376 24452 11395 24508
rect 11301 24428 11395 24452
rect 11301 24372 11320 24428
rect 11376 24372 11395 24428
rect 11301 24348 11395 24372
rect 11301 24292 11320 24348
rect 11376 24292 11395 24348
rect 11301 24264 11395 24292
rect 14191 24588 14285 24616
rect 14191 24532 14210 24588
rect 14266 24532 14285 24588
rect 14191 24508 14285 24532
rect 14191 24452 14210 24508
rect 14266 24452 14285 24508
rect 14191 24428 14285 24452
rect 14191 24372 14210 24428
rect 14266 24372 14285 24428
rect 14191 24348 14285 24372
rect 14191 24292 14210 24348
rect 14266 24292 14285 24348
rect 14191 24264 14285 24292
rect 17081 24588 17175 24616
rect 17081 24532 17100 24588
rect 17156 24532 17175 24588
rect 17081 24508 17175 24532
rect 17081 24452 17100 24508
rect 17156 24452 17175 24508
rect 17081 24428 17175 24452
rect 17081 24372 17100 24428
rect 17156 24372 17175 24428
rect 17081 24348 17175 24372
rect 17081 24292 17100 24348
rect 17156 24292 17175 24348
rect 17081 24264 17175 24292
rect 19971 24588 20065 24616
rect 19971 24532 19990 24588
rect 20046 24532 20065 24588
rect 19971 24508 20065 24532
rect 19971 24452 19990 24508
rect 20046 24452 20065 24508
rect 19971 24428 20065 24452
rect 19971 24372 19990 24428
rect 20046 24372 20065 24428
rect 19971 24348 20065 24372
rect 19971 24292 19990 24348
rect 20046 24292 20065 24348
rect 19971 24264 20065 24292
rect 22861 24588 22955 24616
rect 22861 24532 22880 24588
rect 22936 24532 22955 24588
rect 22861 24508 22955 24532
rect 22861 24452 22880 24508
rect 22936 24452 22955 24508
rect 22861 24428 22955 24452
rect 22861 24372 22880 24428
rect 22936 24372 22955 24428
rect 22861 24348 22955 24372
rect 22861 24292 22880 24348
rect 22936 24292 22955 24348
rect 22861 24264 22955 24292
rect 25751 24588 25845 24616
rect 25751 24532 25770 24588
rect 25826 24532 25845 24588
rect 25751 24508 25845 24532
rect 25751 24452 25770 24508
rect 25826 24452 25845 24508
rect 25751 24428 25845 24452
rect 25751 24372 25770 24428
rect 25826 24372 25845 24428
rect 25751 24348 25845 24372
rect 25751 24292 25770 24348
rect 25826 24292 25845 24348
rect 25751 24264 25845 24292
rect 28641 24588 28735 24616
rect 28641 24532 28660 24588
rect 28716 24532 28735 24588
rect 28641 24508 28735 24532
rect 28641 24452 28660 24508
rect 28716 24452 28735 24508
rect 28641 24428 28735 24452
rect 28641 24372 28660 24428
rect 28716 24372 28735 24428
rect 28641 24348 28735 24372
rect 28641 24292 28660 24348
rect 28716 24292 28735 24348
rect 28641 24264 28735 24292
rect 31531 24588 31625 24616
rect 31531 24532 31550 24588
rect 31606 24532 31625 24588
rect 31531 24508 31625 24532
rect 31531 24452 31550 24508
rect 31606 24452 31625 24508
rect 31531 24428 31625 24452
rect 31531 24372 31550 24428
rect 31606 24372 31625 24428
rect 31531 24348 31625 24372
rect 31531 24292 31550 24348
rect 31606 24292 31625 24348
rect 31531 24264 31625 24292
rect 34421 24588 34515 24616
rect 34421 24532 34440 24588
rect 34496 24532 34515 24588
rect 34421 24508 34515 24532
rect 34421 24452 34440 24508
rect 34496 24452 34515 24508
rect 34421 24428 34515 24452
rect 34421 24372 34440 24428
rect 34496 24372 34515 24428
rect 34421 24348 34515 24372
rect 34421 24292 34440 24348
rect 34496 24292 34515 24348
rect 34421 24264 34515 24292
rect 37311 24588 37405 24616
rect 37311 24532 37330 24588
rect 37386 24532 37405 24588
rect 37311 24508 37405 24532
rect 37311 24452 37330 24508
rect 37386 24452 37405 24508
rect 37311 24428 37405 24452
rect 37311 24372 37330 24428
rect 37386 24372 37405 24428
rect 37311 24348 37405 24372
rect 37311 24292 37330 24348
rect 37386 24292 37405 24348
rect 37311 24264 37405 24292
rect 40201 24588 40295 24616
rect 40201 24532 40220 24588
rect 40276 24532 40295 24588
rect 40201 24508 40295 24532
rect 40201 24452 40220 24508
rect 40276 24452 40295 24508
rect 40201 24428 40295 24452
rect 40201 24372 40220 24428
rect 40276 24372 40295 24428
rect 40201 24348 40295 24372
rect 40201 24292 40220 24348
rect 40276 24292 40295 24348
rect 40201 24264 40295 24292
rect 43091 24588 43185 24616
rect 43091 24532 43110 24588
rect 43166 24532 43185 24588
rect 43091 24508 43185 24532
rect 43091 24452 43110 24508
rect 43166 24452 43185 24508
rect 43091 24428 43185 24452
rect 43091 24372 43110 24428
rect 43166 24372 43185 24428
rect 43091 24348 43185 24372
rect 43091 24292 43110 24348
rect 43166 24292 43185 24348
rect 43091 24264 43185 24292
rect 45981 24588 46075 24616
rect 45981 24532 46000 24588
rect 46056 24532 46075 24588
rect 45981 24508 46075 24532
rect 45981 24452 46000 24508
rect 46056 24452 46075 24508
rect 45981 24428 46075 24452
rect 45981 24372 46000 24428
rect 46056 24372 46075 24428
rect 45981 24348 46075 24372
rect 45981 24292 46000 24348
rect 46056 24292 46075 24348
rect 45981 24264 46075 24292
rect 48989 24588 49083 24616
rect 48989 24532 49008 24588
rect 49064 24532 49083 24588
rect 48989 24508 49083 24532
rect 48989 24452 49008 24508
rect 49064 24452 49083 24508
rect 48989 24428 49083 24452
rect 48989 24372 49008 24428
rect 49064 24372 49083 24428
rect 48989 24348 49083 24372
rect 48989 24292 49008 24348
rect 49064 24292 49083 24348
rect 48989 24264 49083 24292
rect 52210 24588 52320 24616
rect 52210 24532 52237 24588
rect 52293 24532 52320 24588
rect 52210 24508 52320 24532
rect 52210 24452 52237 24508
rect 52293 24452 52320 24508
rect 52210 24428 52320 24452
rect 52210 24372 52237 24428
rect 52293 24372 52320 24428
rect 52210 24348 52320 24372
rect 52210 24292 52237 24348
rect 52293 24292 52320 24348
rect 52210 24264 52320 24292
rect 53602 24588 53730 24616
rect 53602 24532 53638 24588
rect 53694 24532 53730 24588
rect 53602 24508 53730 24532
rect 53602 24452 53638 24508
rect 53694 24452 53730 24508
rect 53602 24428 53730 24452
rect 53602 24372 53638 24428
rect 53694 24372 53730 24428
rect 53602 24348 53730 24372
rect 53602 24292 53638 24348
rect 53694 24292 53730 24348
rect 53602 24264 53730 24292
rect 53770 24588 53898 24616
rect 53770 24532 53806 24588
rect 53862 24532 53898 24588
rect 53770 24508 53898 24532
rect 53770 24452 53806 24508
rect 53862 24452 53898 24508
rect 53770 24428 53898 24452
rect 53770 24372 53806 24428
rect 53862 24372 53898 24428
rect 53770 24348 53898 24372
rect 53770 24292 53806 24348
rect 53862 24292 53898 24348
rect 53770 24264 53898 24292
rect 54514 24588 54642 24616
rect 54514 24532 54550 24588
rect 54606 24532 54642 24588
rect 54514 24508 54642 24532
rect 54514 24452 54550 24508
rect 54606 24452 54642 24508
rect 54514 24428 54642 24452
rect 54514 24372 54550 24428
rect 54606 24372 54642 24428
rect 54514 24348 54642 24372
rect 54514 24292 54550 24348
rect 54606 24292 54642 24348
rect 54514 24264 54642 24292
rect 54910 24588 55026 24616
rect 54910 24532 54940 24588
rect 54996 24532 55026 24588
rect 54910 24508 55026 24532
rect 54910 24452 54940 24508
rect 54996 24452 55026 24508
rect 54910 24428 55026 24452
rect 54910 24372 54940 24428
rect 54996 24372 55026 24428
rect 54910 24348 55026 24372
rect 54910 24292 54940 24348
rect 54996 24292 55026 24348
rect 54910 24264 55026 24292
rect 55620 24588 55748 24616
rect 55620 24532 55656 24588
rect 55712 24532 55748 24588
rect 55620 24508 55748 24532
rect 55620 24452 55656 24508
rect 55712 24452 55748 24508
rect 55620 24428 55748 24452
rect 55620 24372 55656 24428
rect 55712 24372 55748 24428
rect 55620 24348 55748 24372
rect 55620 24292 55656 24348
rect 55712 24292 55748 24348
rect 55620 24264 55748 24292
rect 56198 24588 56326 24616
rect 56198 24532 56234 24588
rect 56290 24532 56326 24588
rect 56198 24508 56326 24532
rect 56198 24452 56234 24508
rect 56290 24452 56326 24508
rect 56198 24428 56326 24452
rect 56198 24372 56234 24428
rect 56290 24372 56326 24428
rect 56198 24348 56326 24372
rect 56198 24292 56234 24348
rect 56290 24292 56326 24348
rect 56198 24264 56326 24292
rect 56649 24588 56765 24616
rect 56649 24532 56679 24588
rect 56735 24532 56765 24588
rect 56649 24508 56765 24532
rect 56649 24452 56679 24508
rect 56735 24452 56765 24508
rect 56649 24428 56765 24452
rect 56649 24372 56679 24428
rect 56735 24372 56765 24428
rect 56649 24348 56765 24372
rect 56649 24292 56679 24348
rect 56735 24292 56765 24348
rect 56649 24264 56765 24292
rect 56953 24588 57069 24616
rect 56953 24532 56983 24588
rect 57039 24532 57069 24588
rect 56953 24508 57069 24532
rect 56953 24452 56983 24508
rect 57039 24452 57069 24508
rect 56953 24428 57069 24452
rect 56953 24372 56983 24428
rect 57039 24372 57069 24428
rect 56953 24348 57069 24372
rect 56953 24292 56983 24348
rect 57039 24292 57069 24348
rect 56953 24264 57069 24292
rect 57795 24588 57911 24616
rect 57795 24532 57825 24588
rect 57881 24532 57911 24588
rect 57795 24508 57911 24532
rect 57795 24452 57825 24508
rect 57881 24452 57911 24508
rect 57795 24428 57911 24452
rect 57795 24372 57825 24428
rect 57881 24372 57911 24428
rect 57795 24348 57911 24372
rect 57795 24292 57825 24348
rect 57881 24292 57911 24348
rect 57795 24264 57911 24292
rect 58461 24588 58525 24616
rect 58461 24532 58465 24588
rect 58521 24532 58525 24588
rect 58461 24508 58525 24532
rect 58461 24452 58465 24508
rect 58521 24452 58525 24508
rect 58461 24428 58525 24452
rect 58461 24372 58465 24428
rect 58521 24372 58525 24428
rect 58461 24348 58525 24372
rect 58461 24292 58465 24348
rect 58521 24292 58525 24348
rect 58461 24264 58525 24292
rect 59018 24588 59134 24616
rect 59018 24532 59048 24588
rect 59104 24532 59134 24588
rect 59018 24508 59134 24532
rect 59018 24452 59048 24508
rect 59104 24452 59134 24508
rect 59018 24428 59134 24452
rect 59018 24372 59048 24428
rect 59104 24372 59134 24428
rect 59018 24348 59134 24372
rect 59018 24292 59048 24348
rect 59104 24292 59134 24348
rect 59018 24264 59134 24292
rect 60296 24588 60412 24616
rect 60296 24532 60326 24588
rect 60382 24532 60412 24588
rect 60296 24508 60412 24532
rect 60296 24452 60326 24508
rect 60382 24452 60412 24508
rect 60296 24428 60412 24452
rect 60296 24372 60326 24428
rect 60382 24372 60412 24428
rect 60296 24348 60412 24372
rect 60296 24292 60326 24348
rect 60382 24292 60412 24348
rect 60296 24264 60412 24292
rect 60454 24588 60570 24616
rect 60454 24532 60484 24588
rect 60540 24532 60570 24588
rect 60454 24508 60570 24532
rect 60454 24452 60484 24508
rect 60540 24452 60570 24508
rect 60454 24428 60570 24452
rect 60454 24372 60484 24428
rect 60540 24372 60570 24428
rect 60454 24348 60570 24372
rect 60454 24292 60484 24348
rect 60540 24292 60570 24348
rect 60454 24264 60570 24292
rect 62509 24588 62683 24616
rect 62509 24532 62528 24588
rect 62584 24532 62608 24588
rect 62664 24532 62683 24588
rect 62509 24508 62683 24532
rect 62509 24452 62528 24508
rect 62584 24452 62608 24508
rect 62664 24452 62683 24508
rect 62509 24428 62683 24452
rect 62509 24372 62528 24428
rect 62584 24372 62608 24428
rect 62664 24372 62683 24428
rect 62509 24348 62683 24372
rect 62509 24292 62528 24348
rect 62584 24292 62608 24348
rect 62664 24292 62683 24348
rect 62509 24264 62683 24292
rect 2152 22236 2352 22264
rect 2152 22180 2184 22236
rect 2240 22180 2264 22236
rect 2320 22180 2352 22236
rect 2152 22156 2352 22180
rect 2152 22100 2184 22156
rect 2240 22100 2264 22156
rect 2320 22100 2352 22156
rect 2152 22076 2352 22100
rect 2152 22020 2184 22076
rect 2240 22020 2264 22076
rect 2320 22020 2352 22076
rect 2152 21996 2352 22020
rect 2152 21940 2184 21996
rect 2240 21940 2264 21996
rect 2320 21940 2352 21996
rect 2152 21912 2352 21940
rect 5374 22236 5468 22264
rect 5374 22180 5393 22236
rect 5449 22180 5468 22236
rect 5374 22156 5468 22180
rect 5374 22100 5393 22156
rect 5449 22100 5468 22156
rect 5374 22076 5468 22100
rect 5374 22020 5393 22076
rect 5449 22020 5468 22076
rect 5374 21996 5468 22020
rect 5374 21940 5393 21996
rect 5449 21940 5468 21996
rect 5374 21912 5468 21940
rect 8264 22236 8358 22264
rect 8264 22180 8283 22236
rect 8339 22180 8358 22236
rect 8264 22156 8358 22180
rect 8264 22100 8283 22156
rect 8339 22100 8358 22156
rect 8264 22076 8358 22100
rect 8264 22020 8283 22076
rect 8339 22020 8358 22076
rect 8264 21996 8358 22020
rect 8264 21940 8283 21996
rect 8339 21940 8358 21996
rect 8264 21912 8358 21940
rect 11154 22236 11248 22264
rect 11154 22180 11173 22236
rect 11229 22180 11248 22236
rect 11154 22156 11248 22180
rect 11154 22100 11173 22156
rect 11229 22100 11248 22156
rect 11154 22076 11248 22100
rect 11154 22020 11173 22076
rect 11229 22020 11248 22076
rect 11154 21996 11248 22020
rect 11154 21940 11173 21996
rect 11229 21940 11248 21996
rect 11154 21912 11248 21940
rect 14044 22236 14138 22264
rect 14044 22180 14063 22236
rect 14119 22180 14138 22236
rect 14044 22156 14138 22180
rect 14044 22100 14063 22156
rect 14119 22100 14138 22156
rect 14044 22076 14138 22100
rect 14044 22020 14063 22076
rect 14119 22020 14138 22076
rect 14044 21996 14138 22020
rect 14044 21940 14063 21996
rect 14119 21940 14138 21996
rect 14044 21912 14138 21940
rect 16934 22236 17028 22264
rect 16934 22180 16953 22236
rect 17009 22180 17028 22236
rect 16934 22156 17028 22180
rect 16934 22100 16953 22156
rect 17009 22100 17028 22156
rect 16934 22076 17028 22100
rect 16934 22020 16953 22076
rect 17009 22020 17028 22076
rect 16934 21996 17028 22020
rect 16934 21940 16953 21996
rect 17009 21940 17028 21996
rect 16934 21912 17028 21940
rect 19824 22236 19918 22264
rect 19824 22180 19843 22236
rect 19899 22180 19918 22236
rect 19824 22156 19918 22180
rect 19824 22100 19843 22156
rect 19899 22100 19918 22156
rect 19824 22076 19918 22100
rect 19824 22020 19843 22076
rect 19899 22020 19918 22076
rect 19824 21996 19918 22020
rect 19824 21940 19843 21996
rect 19899 21940 19918 21996
rect 19824 21912 19918 21940
rect 22714 22236 22808 22264
rect 22714 22180 22733 22236
rect 22789 22180 22808 22236
rect 22714 22156 22808 22180
rect 22714 22100 22733 22156
rect 22789 22100 22808 22156
rect 22714 22076 22808 22100
rect 22714 22020 22733 22076
rect 22789 22020 22808 22076
rect 22714 21996 22808 22020
rect 22714 21940 22733 21996
rect 22789 21940 22808 21996
rect 22714 21912 22808 21940
rect 25604 22236 25698 22264
rect 25604 22180 25623 22236
rect 25679 22180 25698 22236
rect 25604 22156 25698 22180
rect 25604 22100 25623 22156
rect 25679 22100 25698 22156
rect 25604 22076 25698 22100
rect 25604 22020 25623 22076
rect 25679 22020 25698 22076
rect 25604 21996 25698 22020
rect 25604 21940 25623 21996
rect 25679 21940 25698 21996
rect 25604 21912 25698 21940
rect 28494 22236 28588 22264
rect 28494 22180 28513 22236
rect 28569 22180 28588 22236
rect 28494 22156 28588 22180
rect 28494 22100 28513 22156
rect 28569 22100 28588 22156
rect 28494 22076 28588 22100
rect 28494 22020 28513 22076
rect 28569 22020 28588 22076
rect 28494 21996 28588 22020
rect 28494 21940 28513 21996
rect 28569 21940 28588 21996
rect 28494 21912 28588 21940
rect 31384 22236 31478 22264
rect 31384 22180 31403 22236
rect 31459 22180 31478 22236
rect 31384 22156 31478 22180
rect 31384 22100 31403 22156
rect 31459 22100 31478 22156
rect 31384 22076 31478 22100
rect 31384 22020 31403 22076
rect 31459 22020 31478 22076
rect 31384 21996 31478 22020
rect 31384 21940 31403 21996
rect 31459 21940 31478 21996
rect 31384 21912 31478 21940
rect 34274 22236 34368 22264
rect 34274 22180 34293 22236
rect 34349 22180 34368 22236
rect 34274 22156 34368 22180
rect 34274 22100 34293 22156
rect 34349 22100 34368 22156
rect 34274 22076 34368 22100
rect 34274 22020 34293 22076
rect 34349 22020 34368 22076
rect 34274 21996 34368 22020
rect 34274 21940 34293 21996
rect 34349 21940 34368 21996
rect 34274 21912 34368 21940
rect 37164 22236 37258 22264
rect 37164 22180 37183 22236
rect 37239 22180 37258 22236
rect 37164 22156 37258 22180
rect 37164 22100 37183 22156
rect 37239 22100 37258 22156
rect 37164 22076 37258 22100
rect 37164 22020 37183 22076
rect 37239 22020 37258 22076
rect 37164 21996 37258 22020
rect 37164 21940 37183 21996
rect 37239 21940 37258 21996
rect 37164 21912 37258 21940
rect 40054 22236 40148 22264
rect 40054 22180 40073 22236
rect 40129 22180 40148 22236
rect 40054 22156 40148 22180
rect 40054 22100 40073 22156
rect 40129 22100 40148 22156
rect 40054 22076 40148 22100
rect 40054 22020 40073 22076
rect 40129 22020 40148 22076
rect 40054 21996 40148 22020
rect 40054 21940 40073 21996
rect 40129 21940 40148 21996
rect 40054 21912 40148 21940
rect 42944 22236 43038 22264
rect 42944 22180 42963 22236
rect 43019 22180 43038 22236
rect 42944 22156 43038 22180
rect 42944 22100 42963 22156
rect 43019 22100 43038 22156
rect 42944 22076 43038 22100
rect 42944 22020 42963 22076
rect 43019 22020 43038 22076
rect 42944 21996 43038 22020
rect 42944 21940 42963 21996
rect 43019 21940 43038 21996
rect 42944 21912 43038 21940
rect 45834 22236 45928 22264
rect 45834 22180 45853 22236
rect 45909 22180 45928 22236
rect 45834 22156 45928 22180
rect 45834 22100 45853 22156
rect 45909 22100 45928 22156
rect 45834 22076 45928 22100
rect 45834 22020 45853 22076
rect 45909 22020 45928 22076
rect 45834 21996 45928 22020
rect 45834 21940 45853 21996
rect 45909 21940 45928 21996
rect 45834 21912 45928 21940
rect 48781 22236 48875 22264
rect 48781 22180 48800 22236
rect 48856 22180 48875 22236
rect 48781 22156 48875 22180
rect 48781 22100 48800 22156
rect 48856 22100 48875 22156
rect 48781 22076 48875 22100
rect 48781 22020 48800 22076
rect 48856 22020 48875 22076
rect 48781 21996 48875 22020
rect 48781 21940 48800 21996
rect 48856 21940 48875 21996
rect 48781 21912 48875 21940
rect 49630 22236 49830 22264
rect 49630 22180 49662 22236
rect 49718 22180 49742 22236
rect 49798 22180 49830 22236
rect 49630 22156 49830 22180
rect 49630 22100 49662 22156
rect 49718 22100 49742 22156
rect 49798 22100 49830 22156
rect 49630 22076 49830 22100
rect 49630 22020 49662 22076
rect 49718 22020 49742 22076
rect 49798 22020 49830 22076
rect 49630 21996 49830 22020
rect 49630 21940 49662 21996
rect 49718 21940 49742 21996
rect 49798 21940 49830 21996
rect 49630 21912 49830 21940
rect 52920 22236 53048 22264
rect 52920 22180 52956 22236
rect 53012 22180 53048 22236
rect 52920 22156 53048 22180
rect 52920 22100 52956 22156
rect 53012 22100 53048 22156
rect 52920 22076 53048 22100
rect 52920 22020 52956 22076
rect 53012 22020 53048 22076
rect 52920 21996 53048 22020
rect 52920 21940 52956 21996
rect 53012 21940 53048 21996
rect 52920 21912 53048 21940
rect 53078 22236 53206 22264
rect 53078 22180 53114 22236
rect 53170 22180 53206 22236
rect 53078 22156 53206 22180
rect 53078 22100 53114 22156
rect 53170 22100 53206 22156
rect 53078 22076 53206 22100
rect 53078 22020 53114 22076
rect 53170 22020 53206 22076
rect 53078 21996 53206 22020
rect 53078 21940 53114 21996
rect 53170 21940 53206 21996
rect 53078 21912 53206 21940
rect 53434 22236 53562 22264
rect 53434 22180 53470 22236
rect 53526 22180 53562 22236
rect 53434 22156 53562 22180
rect 53434 22100 53470 22156
rect 53526 22100 53562 22156
rect 53434 22076 53562 22100
rect 53434 22020 53470 22076
rect 53526 22020 53562 22076
rect 53434 21996 53562 22020
rect 53434 21940 53470 21996
rect 53526 21940 53562 21996
rect 53434 21912 53562 21940
rect 54752 22236 54880 22264
rect 54752 22180 54788 22236
rect 54844 22180 54880 22236
rect 54752 22156 54880 22180
rect 54752 22100 54788 22156
rect 54844 22100 54880 22156
rect 54752 22076 54880 22100
rect 54752 22020 54788 22076
rect 54844 22020 54880 22076
rect 54752 21996 54880 22020
rect 54752 21940 54788 21996
rect 54844 21940 54880 21996
rect 54752 21912 54880 21940
rect 55345 22236 55473 22264
rect 55345 22180 55381 22236
rect 55437 22180 55473 22236
rect 55345 22156 55473 22180
rect 55345 22100 55381 22156
rect 55437 22100 55473 22156
rect 55345 22076 55473 22100
rect 55345 22020 55381 22076
rect 55437 22020 55473 22076
rect 55345 21996 55473 22020
rect 55345 21940 55381 21996
rect 55437 21940 55473 21996
rect 55345 21912 55473 21940
rect 56491 22236 56619 22264
rect 56491 22180 56527 22236
rect 56583 22180 56619 22236
rect 56491 22156 56619 22180
rect 56491 22100 56527 22156
rect 56583 22100 56619 22156
rect 56491 22076 56619 22100
rect 56491 22020 56527 22076
rect 56583 22020 56619 22076
rect 56491 21996 56619 22020
rect 56491 21940 56527 21996
rect 56583 21940 56619 21996
rect 56491 21912 56619 21940
rect 57941 22236 58121 22264
rect 57941 22180 57963 22236
rect 58019 22180 58043 22236
rect 58099 22180 58121 22236
rect 57941 22156 58121 22180
rect 57941 22100 57963 22156
rect 58019 22100 58043 22156
rect 58099 22100 58121 22156
rect 57941 22076 58121 22100
rect 57941 22020 57963 22076
rect 58019 22020 58043 22076
rect 58099 22020 58121 22076
rect 57941 21996 58121 22020
rect 57941 21940 57963 21996
rect 58019 21940 58043 21996
rect 58099 21940 58121 21996
rect 57941 21912 58121 21940
rect 59164 22236 59304 22264
rect 59164 22180 59206 22236
rect 59262 22180 59304 22236
rect 59164 22156 59304 22180
rect 59164 22100 59206 22156
rect 59262 22100 59304 22156
rect 59164 22076 59304 22100
rect 59164 22020 59206 22076
rect 59262 22020 59304 22076
rect 59164 21996 59304 22020
rect 59164 21940 59206 21996
rect 59262 21940 59304 21996
rect 59164 21912 59304 21940
rect 59334 22236 59450 22264
rect 59334 22180 59364 22236
rect 59420 22180 59450 22236
rect 59334 22156 59450 22180
rect 59334 22100 59364 22156
rect 59420 22100 59450 22156
rect 59334 22076 59450 22100
rect 59334 22020 59364 22076
rect 59420 22020 59450 22076
rect 59334 21996 59450 22020
rect 59334 21940 59364 21996
rect 59420 21940 59450 21996
rect 59334 21912 59450 21940
rect 59642 22236 59758 22264
rect 59642 22180 59672 22236
rect 59728 22180 59758 22236
rect 59642 22156 59758 22180
rect 59642 22100 59672 22156
rect 59728 22100 59758 22156
rect 59642 22076 59758 22100
rect 59642 22020 59672 22076
rect 59728 22020 59758 22076
rect 59642 21996 59758 22020
rect 59642 21940 59672 21996
rect 59728 21940 59758 21996
rect 59642 21912 59758 21940
rect 59788 22236 59904 22264
rect 59788 22180 59818 22236
rect 59874 22180 59904 22236
rect 59788 22156 59904 22180
rect 59788 22100 59818 22156
rect 59874 22100 59904 22156
rect 59788 22076 59904 22100
rect 59788 22020 59818 22076
rect 59874 22020 59904 22076
rect 59788 21996 59904 22020
rect 59788 21940 59818 21996
rect 59874 21940 59904 21996
rect 59788 21912 59904 21940
rect 59934 22236 60110 22264
rect 59934 22180 59954 22236
rect 60010 22180 60034 22236
rect 60090 22180 60110 22236
rect 59934 22156 60110 22180
rect 59934 22100 59954 22156
rect 60010 22100 60034 22156
rect 60090 22100 60110 22156
rect 59934 22076 60110 22100
rect 59934 22020 59954 22076
rect 60010 22020 60034 22076
rect 60090 22020 60110 22076
rect 59934 21996 60110 22020
rect 59934 21940 59954 21996
rect 60010 21940 60034 21996
rect 60090 21940 60110 21996
rect 59934 21912 60110 21940
rect 62307 22236 62481 22264
rect 62307 22180 62326 22236
rect 62382 22180 62406 22236
rect 62462 22180 62481 22236
rect 62307 22156 62481 22180
rect 62307 22100 62326 22156
rect 62382 22100 62406 22156
rect 62462 22100 62481 22156
rect 62307 22076 62481 22100
rect 62307 22020 62326 22076
rect 62382 22020 62406 22076
rect 62462 22020 62481 22076
rect 62307 21996 62481 22020
rect 62307 21940 62326 21996
rect 62382 21940 62406 21996
rect 62462 21940 62481 21996
rect 62307 21912 62481 21940
rect 2020 14588 2124 14616
rect 2020 14532 2044 14588
rect 2100 14532 2124 14588
rect 2020 14508 2124 14532
rect 2020 14452 2044 14508
rect 2100 14452 2124 14508
rect 2020 14428 2124 14452
rect 2020 14372 2044 14428
rect 2100 14372 2124 14428
rect 2020 14348 2124 14372
rect 2020 14292 2044 14348
rect 2100 14292 2124 14348
rect 2020 14264 2124 14292
rect 5521 14588 5615 14616
rect 5521 14532 5540 14588
rect 5596 14532 5615 14588
rect 5521 14508 5615 14532
rect 5521 14452 5540 14508
rect 5596 14452 5615 14508
rect 5521 14428 5615 14452
rect 5521 14372 5540 14428
rect 5596 14372 5615 14428
rect 5521 14348 5615 14372
rect 5521 14292 5540 14348
rect 5596 14292 5615 14348
rect 5521 14264 5615 14292
rect 8411 14588 8505 14616
rect 8411 14532 8430 14588
rect 8486 14532 8505 14588
rect 8411 14508 8505 14532
rect 8411 14452 8430 14508
rect 8486 14452 8505 14508
rect 8411 14428 8505 14452
rect 8411 14372 8430 14428
rect 8486 14372 8505 14428
rect 8411 14348 8505 14372
rect 8411 14292 8430 14348
rect 8486 14292 8505 14348
rect 8411 14264 8505 14292
rect 11301 14588 11395 14616
rect 11301 14532 11320 14588
rect 11376 14532 11395 14588
rect 11301 14508 11395 14532
rect 11301 14452 11320 14508
rect 11376 14452 11395 14508
rect 11301 14428 11395 14452
rect 11301 14372 11320 14428
rect 11376 14372 11395 14428
rect 11301 14348 11395 14372
rect 11301 14292 11320 14348
rect 11376 14292 11395 14348
rect 11301 14264 11395 14292
rect 14191 14588 14285 14616
rect 14191 14532 14210 14588
rect 14266 14532 14285 14588
rect 14191 14508 14285 14532
rect 14191 14452 14210 14508
rect 14266 14452 14285 14508
rect 14191 14428 14285 14452
rect 14191 14372 14210 14428
rect 14266 14372 14285 14428
rect 14191 14348 14285 14372
rect 14191 14292 14210 14348
rect 14266 14292 14285 14348
rect 14191 14264 14285 14292
rect 17081 14588 17175 14616
rect 17081 14532 17100 14588
rect 17156 14532 17175 14588
rect 17081 14508 17175 14532
rect 17081 14452 17100 14508
rect 17156 14452 17175 14508
rect 17081 14428 17175 14452
rect 17081 14372 17100 14428
rect 17156 14372 17175 14428
rect 17081 14348 17175 14372
rect 17081 14292 17100 14348
rect 17156 14292 17175 14348
rect 17081 14264 17175 14292
rect 19971 14588 20065 14616
rect 19971 14532 19990 14588
rect 20046 14532 20065 14588
rect 19971 14508 20065 14532
rect 19971 14452 19990 14508
rect 20046 14452 20065 14508
rect 19971 14428 20065 14452
rect 19971 14372 19990 14428
rect 20046 14372 20065 14428
rect 19971 14348 20065 14372
rect 19971 14292 19990 14348
rect 20046 14292 20065 14348
rect 19971 14264 20065 14292
rect 22861 14588 22955 14616
rect 22861 14532 22880 14588
rect 22936 14532 22955 14588
rect 22861 14508 22955 14532
rect 22861 14452 22880 14508
rect 22936 14452 22955 14508
rect 22861 14428 22955 14452
rect 22861 14372 22880 14428
rect 22936 14372 22955 14428
rect 22861 14348 22955 14372
rect 22861 14292 22880 14348
rect 22936 14292 22955 14348
rect 22861 14264 22955 14292
rect 25751 14588 25845 14616
rect 25751 14532 25770 14588
rect 25826 14532 25845 14588
rect 25751 14508 25845 14532
rect 25751 14452 25770 14508
rect 25826 14452 25845 14508
rect 25751 14428 25845 14452
rect 25751 14372 25770 14428
rect 25826 14372 25845 14428
rect 25751 14348 25845 14372
rect 25751 14292 25770 14348
rect 25826 14292 25845 14348
rect 25751 14264 25845 14292
rect 28641 14588 28735 14616
rect 28641 14532 28660 14588
rect 28716 14532 28735 14588
rect 28641 14508 28735 14532
rect 28641 14452 28660 14508
rect 28716 14452 28735 14508
rect 28641 14428 28735 14452
rect 28641 14372 28660 14428
rect 28716 14372 28735 14428
rect 28641 14348 28735 14372
rect 28641 14292 28660 14348
rect 28716 14292 28735 14348
rect 28641 14264 28735 14292
rect 31531 14588 31625 14616
rect 31531 14532 31550 14588
rect 31606 14532 31625 14588
rect 31531 14508 31625 14532
rect 31531 14452 31550 14508
rect 31606 14452 31625 14508
rect 31531 14428 31625 14452
rect 31531 14372 31550 14428
rect 31606 14372 31625 14428
rect 31531 14348 31625 14372
rect 31531 14292 31550 14348
rect 31606 14292 31625 14348
rect 31531 14264 31625 14292
rect 34421 14588 34515 14616
rect 34421 14532 34440 14588
rect 34496 14532 34515 14588
rect 34421 14508 34515 14532
rect 34421 14452 34440 14508
rect 34496 14452 34515 14508
rect 34421 14428 34515 14452
rect 34421 14372 34440 14428
rect 34496 14372 34515 14428
rect 34421 14348 34515 14372
rect 34421 14292 34440 14348
rect 34496 14292 34515 14348
rect 34421 14264 34515 14292
rect 37311 14588 37405 14616
rect 37311 14532 37330 14588
rect 37386 14532 37405 14588
rect 37311 14508 37405 14532
rect 37311 14452 37330 14508
rect 37386 14452 37405 14508
rect 37311 14428 37405 14452
rect 37311 14372 37330 14428
rect 37386 14372 37405 14428
rect 37311 14348 37405 14372
rect 37311 14292 37330 14348
rect 37386 14292 37405 14348
rect 37311 14264 37405 14292
rect 40201 14588 40295 14616
rect 40201 14532 40220 14588
rect 40276 14532 40295 14588
rect 40201 14508 40295 14532
rect 40201 14452 40220 14508
rect 40276 14452 40295 14508
rect 40201 14428 40295 14452
rect 40201 14372 40220 14428
rect 40276 14372 40295 14428
rect 40201 14348 40295 14372
rect 40201 14292 40220 14348
rect 40276 14292 40295 14348
rect 40201 14264 40295 14292
rect 43091 14588 43185 14616
rect 43091 14532 43110 14588
rect 43166 14532 43185 14588
rect 43091 14508 43185 14532
rect 43091 14452 43110 14508
rect 43166 14452 43185 14508
rect 43091 14428 43185 14452
rect 43091 14372 43110 14428
rect 43166 14372 43185 14428
rect 43091 14348 43185 14372
rect 43091 14292 43110 14348
rect 43166 14292 43185 14348
rect 43091 14264 43185 14292
rect 45981 14588 46075 14616
rect 45981 14532 46000 14588
rect 46056 14532 46075 14588
rect 45981 14508 46075 14532
rect 45981 14452 46000 14508
rect 46056 14452 46075 14508
rect 45981 14428 46075 14452
rect 45981 14372 46000 14428
rect 46056 14372 46075 14428
rect 45981 14348 46075 14372
rect 45981 14292 46000 14348
rect 46056 14292 46075 14348
rect 45981 14264 46075 14292
rect 48989 14588 49083 14616
rect 48989 14532 49008 14588
rect 49064 14532 49083 14588
rect 48989 14508 49083 14532
rect 48989 14452 49008 14508
rect 49064 14452 49083 14508
rect 48989 14428 49083 14452
rect 48989 14372 49008 14428
rect 49064 14372 49083 14428
rect 48989 14348 49083 14372
rect 48989 14292 49008 14348
rect 49064 14292 49083 14348
rect 48989 14264 49083 14292
rect 52210 14588 52320 14616
rect 52210 14532 52237 14588
rect 52293 14532 52320 14588
rect 52210 14508 52320 14532
rect 52210 14452 52237 14508
rect 52293 14452 52320 14508
rect 52210 14428 52320 14452
rect 52210 14372 52237 14428
rect 52293 14372 52320 14428
rect 52210 14348 52320 14372
rect 52210 14292 52237 14348
rect 52293 14292 52320 14348
rect 52210 14264 52320 14292
rect 53602 14588 53730 14616
rect 53602 14532 53638 14588
rect 53694 14532 53730 14588
rect 53602 14508 53730 14532
rect 53602 14452 53638 14508
rect 53694 14452 53730 14508
rect 53602 14428 53730 14452
rect 53602 14372 53638 14428
rect 53694 14372 53730 14428
rect 53602 14348 53730 14372
rect 53602 14292 53638 14348
rect 53694 14292 53730 14348
rect 53602 14264 53730 14292
rect 53770 14588 53898 14616
rect 53770 14532 53806 14588
rect 53862 14532 53898 14588
rect 53770 14508 53898 14532
rect 53770 14452 53806 14508
rect 53862 14452 53898 14508
rect 53770 14428 53898 14452
rect 53770 14372 53806 14428
rect 53862 14372 53898 14428
rect 53770 14348 53898 14372
rect 53770 14292 53806 14348
rect 53862 14292 53898 14348
rect 53770 14264 53898 14292
rect 54514 14588 54642 14616
rect 54514 14532 54550 14588
rect 54606 14532 54642 14588
rect 54514 14508 54642 14532
rect 54514 14452 54550 14508
rect 54606 14452 54642 14508
rect 54514 14428 54642 14452
rect 54514 14372 54550 14428
rect 54606 14372 54642 14428
rect 54514 14348 54642 14372
rect 54514 14292 54550 14348
rect 54606 14292 54642 14348
rect 54514 14264 54642 14292
rect 54910 14588 55026 14616
rect 54910 14532 54940 14588
rect 54996 14532 55026 14588
rect 54910 14508 55026 14532
rect 54910 14452 54940 14508
rect 54996 14452 55026 14508
rect 54910 14428 55026 14452
rect 54910 14372 54940 14428
rect 54996 14372 55026 14428
rect 54910 14348 55026 14372
rect 54910 14292 54940 14348
rect 54996 14292 55026 14348
rect 54910 14264 55026 14292
rect 55620 14588 55748 14616
rect 55620 14532 55656 14588
rect 55712 14532 55748 14588
rect 55620 14508 55748 14532
rect 55620 14452 55656 14508
rect 55712 14452 55748 14508
rect 55620 14428 55748 14452
rect 55620 14372 55656 14428
rect 55712 14372 55748 14428
rect 55620 14348 55748 14372
rect 55620 14292 55656 14348
rect 55712 14292 55748 14348
rect 55620 14264 55748 14292
rect 56198 14588 56326 14616
rect 56198 14532 56234 14588
rect 56290 14532 56326 14588
rect 56198 14508 56326 14532
rect 56198 14452 56234 14508
rect 56290 14452 56326 14508
rect 56198 14428 56326 14452
rect 56198 14372 56234 14428
rect 56290 14372 56326 14428
rect 56198 14348 56326 14372
rect 56198 14292 56234 14348
rect 56290 14292 56326 14348
rect 56198 14264 56326 14292
rect 56649 14588 56765 14616
rect 56649 14532 56679 14588
rect 56735 14532 56765 14588
rect 56649 14508 56765 14532
rect 56649 14452 56679 14508
rect 56735 14452 56765 14508
rect 56649 14428 56765 14452
rect 56649 14372 56679 14428
rect 56735 14372 56765 14428
rect 56649 14348 56765 14372
rect 56649 14292 56679 14348
rect 56735 14292 56765 14348
rect 56649 14264 56765 14292
rect 56953 14588 57069 14616
rect 56953 14532 56983 14588
rect 57039 14532 57069 14588
rect 56953 14508 57069 14532
rect 56953 14452 56983 14508
rect 57039 14452 57069 14508
rect 56953 14428 57069 14452
rect 56953 14372 56983 14428
rect 57039 14372 57069 14428
rect 56953 14348 57069 14372
rect 56953 14292 56983 14348
rect 57039 14292 57069 14348
rect 56953 14264 57069 14292
rect 57795 14588 57911 14616
rect 57795 14532 57825 14588
rect 57881 14532 57911 14588
rect 57795 14508 57911 14532
rect 57795 14452 57825 14508
rect 57881 14452 57911 14508
rect 57795 14428 57911 14452
rect 57795 14372 57825 14428
rect 57881 14372 57911 14428
rect 57795 14348 57911 14372
rect 57795 14292 57825 14348
rect 57881 14292 57911 14348
rect 57795 14264 57911 14292
rect 58461 14588 58525 14616
rect 58461 14532 58465 14588
rect 58521 14532 58525 14588
rect 58461 14508 58525 14532
rect 58461 14452 58465 14508
rect 58521 14452 58525 14508
rect 58461 14428 58525 14452
rect 58461 14372 58465 14428
rect 58521 14372 58525 14428
rect 58461 14348 58525 14372
rect 58461 14292 58465 14348
rect 58521 14292 58525 14348
rect 58461 14264 58525 14292
rect 59018 14588 59134 14616
rect 59018 14532 59048 14588
rect 59104 14532 59134 14588
rect 59018 14508 59134 14532
rect 59018 14452 59048 14508
rect 59104 14452 59134 14508
rect 59018 14428 59134 14452
rect 59018 14372 59048 14428
rect 59104 14372 59134 14428
rect 59018 14348 59134 14372
rect 59018 14292 59048 14348
rect 59104 14292 59134 14348
rect 59018 14264 59134 14292
rect 60296 14588 60412 14616
rect 60296 14532 60326 14588
rect 60382 14532 60412 14588
rect 60296 14508 60412 14532
rect 60296 14452 60326 14508
rect 60382 14452 60412 14508
rect 60296 14428 60412 14452
rect 60296 14372 60326 14428
rect 60382 14372 60412 14428
rect 60296 14348 60412 14372
rect 60296 14292 60326 14348
rect 60382 14292 60412 14348
rect 60296 14264 60412 14292
rect 60454 14588 60570 14616
rect 60454 14532 60484 14588
rect 60540 14532 60570 14588
rect 60454 14508 60570 14532
rect 60454 14452 60484 14508
rect 60540 14452 60570 14508
rect 60454 14428 60570 14452
rect 60454 14372 60484 14428
rect 60540 14372 60570 14428
rect 60454 14348 60570 14372
rect 60454 14292 60484 14348
rect 60540 14292 60570 14348
rect 60454 14264 60570 14292
rect 62509 14588 62683 14616
rect 62509 14532 62528 14588
rect 62584 14532 62608 14588
rect 62664 14532 62683 14588
rect 62509 14508 62683 14532
rect 62509 14452 62528 14508
rect 62584 14452 62608 14508
rect 62664 14452 62683 14508
rect 62509 14428 62683 14452
rect 62509 14372 62528 14428
rect 62584 14372 62608 14428
rect 62664 14372 62683 14428
rect 62509 14348 62683 14372
rect 62509 14292 62528 14348
rect 62584 14292 62608 14348
rect 62664 14292 62683 14348
rect 62509 14264 62683 14292
rect 2152 12236 2352 12264
rect 2152 12180 2184 12236
rect 2240 12180 2264 12236
rect 2320 12180 2352 12236
rect 2152 12156 2352 12180
rect 2152 12100 2184 12156
rect 2240 12100 2264 12156
rect 2320 12100 2352 12156
rect 2152 12076 2352 12100
rect 2152 12020 2184 12076
rect 2240 12020 2264 12076
rect 2320 12020 2352 12076
rect 2152 11996 2352 12020
rect 2152 11940 2184 11996
rect 2240 11940 2264 11996
rect 2320 11940 2352 11996
rect 2152 11912 2352 11940
rect 5374 12236 5468 12264
rect 5374 12180 5393 12236
rect 5449 12180 5468 12236
rect 5374 12156 5468 12180
rect 5374 12100 5393 12156
rect 5449 12100 5468 12156
rect 5374 12076 5468 12100
rect 5374 12020 5393 12076
rect 5449 12020 5468 12076
rect 5374 11996 5468 12020
rect 5374 11940 5393 11996
rect 5449 11940 5468 11996
rect 5374 11912 5468 11940
rect 8264 12236 8358 12264
rect 8264 12180 8283 12236
rect 8339 12180 8358 12236
rect 8264 12156 8358 12180
rect 8264 12100 8283 12156
rect 8339 12100 8358 12156
rect 8264 12076 8358 12100
rect 8264 12020 8283 12076
rect 8339 12020 8358 12076
rect 8264 11996 8358 12020
rect 8264 11940 8283 11996
rect 8339 11940 8358 11996
rect 8264 11912 8358 11940
rect 11154 12236 11248 12264
rect 11154 12180 11173 12236
rect 11229 12180 11248 12236
rect 11154 12156 11248 12180
rect 11154 12100 11173 12156
rect 11229 12100 11248 12156
rect 11154 12076 11248 12100
rect 11154 12020 11173 12076
rect 11229 12020 11248 12076
rect 11154 11996 11248 12020
rect 11154 11940 11173 11996
rect 11229 11940 11248 11996
rect 11154 11912 11248 11940
rect 14044 12236 14138 12264
rect 14044 12180 14063 12236
rect 14119 12180 14138 12236
rect 14044 12156 14138 12180
rect 14044 12100 14063 12156
rect 14119 12100 14138 12156
rect 14044 12076 14138 12100
rect 14044 12020 14063 12076
rect 14119 12020 14138 12076
rect 14044 11996 14138 12020
rect 14044 11940 14063 11996
rect 14119 11940 14138 11996
rect 14044 11912 14138 11940
rect 16934 12236 17028 12264
rect 16934 12180 16953 12236
rect 17009 12180 17028 12236
rect 16934 12156 17028 12180
rect 16934 12100 16953 12156
rect 17009 12100 17028 12156
rect 16934 12076 17028 12100
rect 16934 12020 16953 12076
rect 17009 12020 17028 12076
rect 16934 11996 17028 12020
rect 16934 11940 16953 11996
rect 17009 11940 17028 11996
rect 16934 11912 17028 11940
rect 19824 12236 19918 12264
rect 19824 12180 19843 12236
rect 19899 12180 19918 12236
rect 19824 12156 19918 12180
rect 19824 12100 19843 12156
rect 19899 12100 19918 12156
rect 19824 12076 19918 12100
rect 19824 12020 19843 12076
rect 19899 12020 19918 12076
rect 19824 11996 19918 12020
rect 19824 11940 19843 11996
rect 19899 11940 19918 11996
rect 19824 11912 19918 11940
rect 22714 12236 22808 12264
rect 22714 12180 22733 12236
rect 22789 12180 22808 12236
rect 22714 12156 22808 12180
rect 22714 12100 22733 12156
rect 22789 12100 22808 12156
rect 22714 12076 22808 12100
rect 22714 12020 22733 12076
rect 22789 12020 22808 12076
rect 22714 11996 22808 12020
rect 22714 11940 22733 11996
rect 22789 11940 22808 11996
rect 22714 11912 22808 11940
rect 25604 12236 25698 12264
rect 25604 12180 25623 12236
rect 25679 12180 25698 12236
rect 25604 12156 25698 12180
rect 25604 12100 25623 12156
rect 25679 12100 25698 12156
rect 25604 12076 25698 12100
rect 25604 12020 25623 12076
rect 25679 12020 25698 12076
rect 25604 11996 25698 12020
rect 25604 11940 25623 11996
rect 25679 11940 25698 11996
rect 25604 11912 25698 11940
rect 28494 12236 28588 12264
rect 28494 12180 28513 12236
rect 28569 12180 28588 12236
rect 28494 12156 28588 12180
rect 28494 12100 28513 12156
rect 28569 12100 28588 12156
rect 28494 12076 28588 12100
rect 28494 12020 28513 12076
rect 28569 12020 28588 12076
rect 28494 11996 28588 12020
rect 28494 11940 28513 11996
rect 28569 11940 28588 11996
rect 28494 11912 28588 11940
rect 31384 12236 31478 12264
rect 31384 12180 31403 12236
rect 31459 12180 31478 12236
rect 31384 12156 31478 12180
rect 31384 12100 31403 12156
rect 31459 12100 31478 12156
rect 31384 12076 31478 12100
rect 31384 12020 31403 12076
rect 31459 12020 31478 12076
rect 31384 11996 31478 12020
rect 31384 11940 31403 11996
rect 31459 11940 31478 11996
rect 31384 11912 31478 11940
rect 34274 12236 34368 12264
rect 34274 12180 34293 12236
rect 34349 12180 34368 12236
rect 34274 12156 34368 12180
rect 34274 12100 34293 12156
rect 34349 12100 34368 12156
rect 34274 12076 34368 12100
rect 34274 12020 34293 12076
rect 34349 12020 34368 12076
rect 34274 11996 34368 12020
rect 34274 11940 34293 11996
rect 34349 11940 34368 11996
rect 34274 11912 34368 11940
rect 37164 12236 37258 12264
rect 37164 12180 37183 12236
rect 37239 12180 37258 12236
rect 37164 12156 37258 12180
rect 37164 12100 37183 12156
rect 37239 12100 37258 12156
rect 37164 12076 37258 12100
rect 37164 12020 37183 12076
rect 37239 12020 37258 12076
rect 37164 11996 37258 12020
rect 37164 11940 37183 11996
rect 37239 11940 37258 11996
rect 37164 11912 37258 11940
rect 40054 12236 40148 12264
rect 40054 12180 40073 12236
rect 40129 12180 40148 12236
rect 40054 12156 40148 12180
rect 40054 12100 40073 12156
rect 40129 12100 40148 12156
rect 40054 12076 40148 12100
rect 40054 12020 40073 12076
rect 40129 12020 40148 12076
rect 40054 11996 40148 12020
rect 40054 11940 40073 11996
rect 40129 11940 40148 11996
rect 40054 11912 40148 11940
rect 42944 12236 43038 12264
rect 42944 12180 42963 12236
rect 43019 12180 43038 12236
rect 42944 12156 43038 12180
rect 42944 12100 42963 12156
rect 43019 12100 43038 12156
rect 42944 12076 43038 12100
rect 42944 12020 42963 12076
rect 43019 12020 43038 12076
rect 42944 11996 43038 12020
rect 42944 11940 42963 11996
rect 43019 11940 43038 11996
rect 42944 11912 43038 11940
rect 45834 12236 45928 12264
rect 45834 12180 45853 12236
rect 45909 12180 45928 12236
rect 45834 12156 45928 12180
rect 45834 12100 45853 12156
rect 45909 12100 45928 12156
rect 45834 12076 45928 12100
rect 45834 12020 45853 12076
rect 45909 12020 45928 12076
rect 45834 11996 45928 12020
rect 45834 11940 45853 11996
rect 45909 11940 45928 11996
rect 45834 11912 45928 11940
rect 48781 12236 48875 12264
rect 48781 12180 48800 12236
rect 48856 12180 48875 12236
rect 48781 12156 48875 12180
rect 48781 12100 48800 12156
rect 48856 12100 48875 12156
rect 48781 12076 48875 12100
rect 48781 12020 48800 12076
rect 48856 12020 48875 12076
rect 48781 11996 48875 12020
rect 48781 11940 48800 11996
rect 48856 11940 48875 11996
rect 48781 11912 48875 11940
rect 49630 12236 49830 12264
rect 49630 12180 49662 12236
rect 49718 12180 49742 12236
rect 49798 12180 49830 12236
rect 49630 12156 49830 12180
rect 49630 12100 49662 12156
rect 49718 12100 49742 12156
rect 49798 12100 49830 12156
rect 49630 12076 49830 12100
rect 49630 12020 49662 12076
rect 49718 12020 49742 12076
rect 49798 12020 49830 12076
rect 49630 11996 49830 12020
rect 49630 11940 49662 11996
rect 49718 11940 49742 11996
rect 49798 11940 49830 11996
rect 49630 11912 49830 11940
rect 52920 12236 53048 12264
rect 52920 12180 52956 12236
rect 53012 12180 53048 12236
rect 52920 12156 53048 12180
rect 52920 12100 52956 12156
rect 53012 12100 53048 12156
rect 52920 12076 53048 12100
rect 52920 12020 52956 12076
rect 53012 12020 53048 12076
rect 52920 11996 53048 12020
rect 52920 11940 52956 11996
rect 53012 11940 53048 11996
rect 52920 11912 53048 11940
rect 53078 12236 53206 12264
rect 53078 12180 53114 12236
rect 53170 12180 53206 12236
rect 53078 12156 53206 12180
rect 53078 12100 53114 12156
rect 53170 12100 53206 12156
rect 53078 12076 53206 12100
rect 53078 12020 53114 12076
rect 53170 12020 53206 12076
rect 53078 11996 53206 12020
rect 53078 11940 53114 11996
rect 53170 11940 53206 11996
rect 53078 11912 53206 11940
rect 53434 12236 53562 12264
rect 53434 12180 53470 12236
rect 53526 12180 53562 12236
rect 53434 12156 53562 12180
rect 53434 12100 53470 12156
rect 53526 12100 53562 12156
rect 53434 12076 53562 12100
rect 53434 12020 53470 12076
rect 53526 12020 53562 12076
rect 53434 11996 53562 12020
rect 53434 11940 53470 11996
rect 53526 11940 53562 11996
rect 53434 11912 53562 11940
rect 54752 12236 54880 12264
rect 54752 12180 54788 12236
rect 54844 12180 54880 12236
rect 54752 12156 54880 12180
rect 54752 12100 54788 12156
rect 54844 12100 54880 12156
rect 54752 12076 54880 12100
rect 54752 12020 54788 12076
rect 54844 12020 54880 12076
rect 54752 11996 54880 12020
rect 54752 11940 54788 11996
rect 54844 11940 54880 11996
rect 54752 11912 54880 11940
rect 55345 12236 55473 12264
rect 55345 12180 55381 12236
rect 55437 12180 55473 12236
rect 55345 12156 55473 12180
rect 55345 12100 55381 12156
rect 55437 12100 55473 12156
rect 55345 12076 55473 12100
rect 55345 12020 55381 12076
rect 55437 12020 55473 12076
rect 55345 11996 55473 12020
rect 55345 11940 55381 11996
rect 55437 11940 55473 11996
rect 55345 11912 55473 11940
rect 56491 12236 56619 12264
rect 56491 12180 56527 12236
rect 56583 12180 56619 12236
rect 56491 12156 56619 12180
rect 56491 12100 56527 12156
rect 56583 12100 56619 12156
rect 56491 12076 56619 12100
rect 56491 12020 56527 12076
rect 56583 12020 56619 12076
rect 56491 11996 56619 12020
rect 56491 11940 56527 11996
rect 56583 11940 56619 11996
rect 56491 11912 56619 11940
rect 57941 12236 58121 12264
rect 57941 12180 57963 12236
rect 58019 12180 58043 12236
rect 58099 12180 58121 12236
rect 57941 12156 58121 12180
rect 57941 12100 57963 12156
rect 58019 12100 58043 12156
rect 58099 12100 58121 12156
rect 57941 12076 58121 12100
rect 57941 12020 57963 12076
rect 58019 12020 58043 12076
rect 58099 12020 58121 12076
rect 57941 11996 58121 12020
rect 57941 11940 57963 11996
rect 58019 11940 58043 11996
rect 58099 11940 58121 11996
rect 57941 11912 58121 11940
rect 59164 12236 59304 12264
rect 59164 12180 59206 12236
rect 59262 12180 59304 12236
rect 59164 12156 59304 12180
rect 59164 12100 59206 12156
rect 59262 12100 59304 12156
rect 59164 12076 59304 12100
rect 59164 12020 59206 12076
rect 59262 12020 59304 12076
rect 59164 11996 59304 12020
rect 59164 11940 59206 11996
rect 59262 11940 59304 11996
rect 59164 11912 59304 11940
rect 59334 12236 59450 12264
rect 59334 12180 59364 12236
rect 59420 12180 59450 12236
rect 59334 12156 59450 12180
rect 59334 12100 59364 12156
rect 59420 12100 59450 12156
rect 59334 12076 59450 12100
rect 59334 12020 59364 12076
rect 59420 12020 59450 12076
rect 59334 11996 59450 12020
rect 59334 11940 59364 11996
rect 59420 11940 59450 11996
rect 59334 11912 59450 11940
rect 59642 12236 59758 12264
rect 59642 12180 59672 12236
rect 59728 12180 59758 12236
rect 59642 12156 59758 12180
rect 59642 12100 59672 12156
rect 59728 12100 59758 12156
rect 59642 12076 59758 12100
rect 59642 12020 59672 12076
rect 59728 12020 59758 12076
rect 59642 11996 59758 12020
rect 59642 11940 59672 11996
rect 59728 11940 59758 11996
rect 59642 11912 59758 11940
rect 59788 12236 59904 12264
rect 59788 12180 59818 12236
rect 59874 12180 59904 12236
rect 59788 12156 59904 12180
rect 59788 12100 59818 12156
rect 59874 12100 59904 12156
rect 59788 12076 59904 12100
rect 59788 12020 59818 12076
rect 59874 12020 59904 12076
rect 59788 11996 59904 12020
rect 59788 11940 59818 11996
rect 59874 11940 59904 11996
rect 59788 11912 59904 11940
rect 59934 12236 60110 12264
rect 59934 12180 59954 12236
rect 60010 12180 60034 12236
rect 60090 12180 60110 12236
rect 59934 12156 60110 12180
rect 59934 12100 59954 12156
rect 60010 12100 60034 12156
rect 60090 12100 60110 12156
rect 59934 12076 60110 12100
rect 59934 12020 59954 12076
rect 60010 12020 60034 12076
rect 60090 12020 60110 12076
rect 59934 11996 60110 12020
rect 59934 11940 59954 11996
rect 60010 11940 60034 11996
rect 60090 11940 60110 11996
rect 59934 11912 60110 11940
rect 62307 12236 62481 12264
rect 62307 12180 62326 12236
rect 62382 12180 62406 12236
rect 62462 12180 62481 12236
rect 62307 12156 62481 12180
rect 62307 12100 62326 12156
rect 62382 12100 62406 12156
rect 62462 12100 62481 12156
rect 62307 12076 62481 12100
rect 62307 12020 62326 12076
rect 62382 12020 62406 12076
rect 62462 12020 62481 12076
rect 62307 11996 62481 12020
rect 62307 11940 62326 11996
rect 62382 11940 62406 11996
rect 62462 11940 62481 11996
rect 62307 11912 62481 11940
rect 63408 10344 63460 10350
rect 63408 10286 63460 10292
rect 59196 7800 59224 8024
rect 59572 7818 59600 8024
rect 61660 7880 61712 7886
rect 61660 7822 61712 7828
rect 59188 7772 59224 7800
rect 59560 7812 59612 7818
rect 52276 7744 52328 7750
rect 30838 7712 30894 7721
rect 52276 7686 52328 7692
rect 30838 7647 30894 7656
rect 30286 7576 30342 7585
rect 30286 7511 30342 7520
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 29090 6760 29146 6769
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 1836 4922 2188 5944
rect 1836 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 2188 4922
rect 1836 3834 2188 4870
rect 1836 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 2188 3834
rect 1836 2746 2188 3782
rect 1836 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 2188 2746
rect 1836 2236 2188 2694
rect 1836 2180 1864 2236
rect 1920 2180 1944 2236
rect 2000 2180 2024 2236
rect 2080 2180 2104 2236
rect 2160 2180 2188 2236
rect 1836 2156 2188 2180
rect 1836 2100 1864 2156
rect 1920 2100 1944 2156
rect 2000 2100 2024 2156
rect 2080 2100 2104 2156
rect 2160 2100 2188 2156
rect 1836 2076 2188 2100
rect 1836 2020 1864 2076
rect 1920 2020 1944 2076
rect 2000 2020 2024 2076
rect 2080 2020 2104 2076
rect 2160 2020 2188 2076
rect 1836 1996 2188 2020
rect 1836 1940 1864 1996
rect 1920 1940 1944 1996
rect 2000 1940 2024 1996
rect 2080 1940 2104 1996
rect 2160 1940 2188 1996
rect 1836 1658 2188 1940
rect 1836 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 2188 1658
rect 1836 1040 2188 1606
rect 4188 5466 4540 5972
rect 4188 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 4540 5466
rect 4188 4588 4540 5414
rect 4188 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4540 4588
rect 4188 4508 4540 4532
rect 4188 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4540 4508
rect 4188 4428 4540 4452
rect 4188 4378 4216 4428
rect 4272 4378 4296 4428
rect 4352 4378 4376 4428
rect 4432 4378 4456 4428
rect 4512 4378 4540 4428
rect 4188 4326 4210 4378
rect 4272 4372 4274 4378
rect 4454 4372 4456 4378
rect 4262 4348 4274 4372
rect 4326 4348 4338 4372
rect 4390 4348 4402 4372
rect 4454 4348 4466 4372
rect 4272 4326 4274 4348
rect 4454 4326 4456 4348
rect 4518 4326 4540 4378
rect 4188 4292 4216 4326
rect 4272 4292 4296 4326
rect 4352 4292 4376 4326
rect 4432 4292 4456 4326
rect 4512 4292 4540 4326
rect 4188 3290 4540 4292
rect 4188 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 4540 3290
rect 4188 2202 4540 3238
rect 4188 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 4540 2202
rect 3148 1284 3200 1290
rect 3148 1226 3200 1232
rect 3160 800 3188 1226
rect 4188 1114 4540 2150
rect 11836 4922 12188 5972
rect 11836 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 12188 4922
rect 11836 3834 12188 4870
rect 11836 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 12188 3834
rect 11836 2746 12188 3782
rect 11836 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 12188 2746
rect 11836 2236 12188 2694
rect 11836 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 12188 2236
rect 11836 2156 12188 2180
rect 11836 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 12188 2156
rect 11836 2076 12188 2100
rect 11836 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 12188 2076
rect 11836 1996 12188 2020
rect 11836 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 12188 1996
rect 11836 1658 12188 1940
rect 11836 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 12188 1658
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 4188 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 4540 1114
rect 4188 1040 4540 1062
rect 5092 1018 5120 1294
rect 11836 1040 12188 1606
rect 14188 5466 14540 5972
rect 14188 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 14540 5466
rect 14188 4588 14540 5414
rect 14188 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 14540 4588
rect 14188 4508 14540 4532
rect 14188 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 14540 4508
rect 14188 4428 14540 4452
rect 14188 4378 14216 4428
rect 14272 4378 14296 4428
rect 14352 4378 14376 4428
rect 14432 4378 14456 4428
rect 14512 4378 14540 4428
rect 14188 4326 14210 4378
rect 14272 4372 14274 4378
rect 14454 4372 14456 4378
rect 14262 4348 14274 4372
rect 14326 4348 14338 4372
rect 14390 4348 14402 4372
rect 14454 4348 14466 4372
rect 14272 4326 14274 4348
rect 14454 4326 14456 4348
rect 14518 4326 14540 4378
rect 14188 4292 14216 4326
rect 14272 4292 14296 4326
rect 14352 4292 14376 4326
rect 14432 4292 14456 4326
rect 14512 4292 14540 4326
rect 14188 3290 14540 4292
rect 21836 4922 22188 5972
rect 23308 5778 23336 6666
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23676 5914 23704 6326
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 24188 5466 24540 5972
rect 24582 5944 24638 5953
rect 24582 5879 24638 5888
rect 24596 5778 24624 5879
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 24780 5710 24808 6598
rect 25872 6588 25924 6594
rect 25872 6530 25924 6536
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24188 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 24540 5466
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 21836 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 22188 4922
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 14738 3360 14794 3369
rect 14738 3295 14794 3304
rect 14188 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 14540 3290
rect 14188 2202 14540 3238
rect 14188 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 14540 2202
rect 14188 1114 14540 2150
rect 14188 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 14540 1114
rect 14188 1040 14540 1062
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 14752 800 14780 3295
rect 17880 3126 17908 3946
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 16396 1964 16448 1970
rect 16396 1906 16448 1912
rect 15292 1352 15344 1358
rect 15292 1294 15344 1300
rect 15304 800 15332 1294
rect 15936 1284 15988 1290
rect 15936 1226 15988 1232
rect 15568 1216 15620 1222
rect 15568 1158 15620 1164
rect 15580 950 15608 1158
rect 15568 944 15620 950
rect 15948 898 15976 1226
rect 15568 886 15620 892
rect 15856 870 15976 898
rect 15856 800 15884 870
rect 16408 800 16436 1906
rect 16960 800 16988 2382
rect 17604 2106 17632 2382
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17592 2100 17644 2106
rect 17592 2042 17644 2048
rect 17788 1358 17816 2246
rect 18248 2106 18276 3470
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18340 2038 18368 2246
rect 18328 2032 18380 2038
rect 18328 1974 18380 1980
rect 18432 1970 18460 2790
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 17500 1352 17552 1358
rect 17500 1294 17552 1300
rect 17776 1352 17828 1358
rect 17776 1294 17828 1300
rect 17512 800 17540 1294
rect 18064 800 18092 1838
rect 18708 1578 18736 2926
rect 18616 1550 18736 1578
rect 18616 800 18644 1550
rect 19076 1358 19104 4082
rect 20272 3738 20300 4082
rect 21836 3834 22188 4870
rect 21836 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 22188 3834
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20548 3194 20576 3470
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 3058 20668 3538
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19168 2650 19196 2926
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19352 1902 19380 2994
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19432 2032 19484 2038
rect 19432 1974 19484 1980
rect 19340 1896 19392 1902
rect 19340 1838 19392 1844
rect 19444 1442 19472 1974
rect 19168 1414 19472 1442
rect 19064 1352 19116 1358
rect 19064 1294 19116 1300
rect 19168 800 19196 1414
rect 19432 1284 19484 1290
rect 19432 1226 19484 1232
rect 19444 882 19472 1226
rect 19432 876 19484 882
rect 19432 818 19484 824
rect 19720 800 19748 2450
rect 19812 1358 19840 2790
rect 19904 2650 19932 2926
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 20272 800 20300 2382
rect 20640 2378 20668 2858
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20732 950 20760 2994
rect 20824 2650 20852 3470
rect 20902 3224 20958 3233
rect 20902 3159 20904 3168
rect 20956 3159 20958 3168
rect 20904 3130 20956 3136
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20720 944 20772 950
rect 20720 886 20772 892
rect 20824 800 20852 2450
rect 20916 2310 20944 3130
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21376 800 21404 2382
rect 21468 2106 21496 2790
rect 21744 2650 21772 2926
rect 21836 2746 22188 3782
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 21836 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 22188 2746
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21744 898 21772 2314
rect 21836 2236 22188 2694
rect 21836 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 22188 2236
rect 21836 2156 22188 2180
rect 21836 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 22188 2156
rect 21836 2076 22188 2100
rect 21836 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 22188 2076
rect 21836 1996 22188 2020
rect 21836 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 22188 1996
rect 21836 1658 22188 1940
rect 21836 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 22188 1658
rect 21836 1040 22188 1606
rect 22296 1290 22324 2858
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22388 1970 22416 2790
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 22284 1284 22336 1290
rect 22284 1226 22336 1232
rect 21744 870 21956 898
rect 21928 800 21956 870
rect 22480 800 22508 3470
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 22848 2922 22876 3062
rect 23124 3058 23152 3334
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23020 2984 23072 2990
rect 23020 2926 23072 2932
rect 22836 2916 22888 2922
rect 22836 2858 22888 2864
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 1358 22600 2790
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22940 1562 22968 2382
rect 22928 1556 22980 1562
rect 22928 1498 22980 1504
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 23032 800 23060 2926
rect 23308 2650 23336 3334
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23204 1896 23256 1902
rect 23492 1850 23520 5034
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23584 3534 23612 3878
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23204 1838 23256 1844
rect 23216 1465 23244 1838
rect 23400 1822 23520 1850
rect 23400 1766 23428 1822
rect 23388 1760 23440 1766
rect 23388 1702 23440 1708
rect 23202 1456 23258 1465
rect 23202 1391 23258 1400
rect 23572 1284 23624 1290
rect 23572 1226 23624 1232
rect 23584 800 23612 1226
rect 23952 1018 23980 5170
rect 24188 4588 24540 5414
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24596 4690 24624 5102
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 24188 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 24540 4588
rect 24188 4508 24540 4532
rect 24188 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 24540 4508
rect 24188 4428 24540 4452
rect 24188 4378 24216 4428
rect 24272 4378 24296 4428
rect 24352 4378 24376 4428
rect 24432 4378 24456 4428
rect 24512 4378 24540 4428
rect 24188 4326 24210 4378
rect 24272 4372 24274 4378
rect 24454 4372 24456 4378
rect 24262 4348 24274 4372
rect 24326 4348 24338 4372
rect 24390 4348 24402 4372
rect 24454 4348 24466 4372
rect 24272 4326 24274 4348
rect 24454 4326 24456 4348
rect 24518 4326 24540 4378
rect 24188 4292 24216 4326
rect 24272 4292 24296 4326
rect 24352 4292 24376 4326
rect 24432 4292 24456 4326
rect 24512 4292 24540 4326
rect 24188 3290 24540 4292
rect 24188 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 24540 3290
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 24044 2650 24072 2926
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23940 1012 23992 1018
rect 23940 954 23992 960
rect 24044 898 24072 2382
rect 24188 2202 24540 3238
rect 24872 3194 24900 5170
rect 24964 3602 24992 6122
rect 25884 5710 25912 6530
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26160 5710 26188 6258
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25976 5370 26004 5646
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25412 5160 25464 5166
rect 26332 5160 26384 5166
rect 25412 5102 25464 5108
rect 25778 5128 25834 5137
rect 25424 4758 25452 5102
rect 26332 5102 26384 5108
rect 25778 5063 25780 5072
rect 25832 5063 25834 5072
rect 25780 5034 25832 5040
rect 26148 5024 26200 5030
rect 26148 4966 26200 4972
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 26160 4486 26188 4966
rect 26252 4826 26280 4966
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 26344 4282 26372 5102
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26712 4554 26740 4966
rect 26700 4548 26752 4554
rect 26700 4490 26752 4496
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24188 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 24540 2202
rect 24188 1114 24540 2150
rect 24596 2106 24624 2382
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 24964 1970 24992 2790
rect 25240 2650 25268 3470
rect 25792 3194 25820 3470
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25884 3233 25912 3402
rect 25870 3224 25926 3233
rect 25780 3188 25832 3194
rect 25870 3159 25926 3168
rect 25780 3130 25832 3136
rect 26068 3126 26096 3674
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26056 3120 26108 3126
rect 26160 3097 26188 3402
rect 26056 3062 26108 3068
rect 26146 3088 26202 3097
rect 26146 3023 26202 3032
rect 26976 3052 27028 3058
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25332 2650 25360 2926
rect 26160 2922 26188 3023
rect 26976 2994 27028 3000
rect 26148 2916 26200 2922
rect 26148 2858 26200 2864
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 24676 1896 24728 1902
rect 24676 1838 24728 1844
rect 24188 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 24540 1114
rect 24188 1040 24540 1062
rect 24044 870 24164 898
rect 24136 800 24164 870
rect 24688 800 24716 1838
rect 25240 800 25268 2382
rect 25884 1970 25912 2518
rect 25976 2514 26004 2790
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 25872 1964 25924 1970
rect 25872 1906 25924 1912
rect 26068 1562 26096 2382
rect 26056 1556 26108 1562
rect 26056 1498 26108 1504
rect 26332 1352 26384 1358
rect 26332 1294 26384 1300
rect 25780 1284 25832 1290
rect 25780 1226 25832 1232
rect 25792 800 25820 1226
rect 26344 800 26372 1294
rect 26528 1222 26556 2790
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 26700 2304 26752 2310
rect 26700 2246 26752 2252
rect 26792 2304 26844 2310
rect 26792 2246 26844 2252
rect 26712 1970 26740 2246
rect 26804 2038 26832 2246
rect 26792 2032 26844 2038
rect 26792 1974 26844 1980
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 26516 1216 26568 1222
rect 26516 1158 26568 1164
rect 26896 800 26924 2382
rect 26988 2106 27016 2994
rect 27080 2990 27108 6190
rect 27158 5264 27214 5273
rect 27158 5199 27214 5208
rect 27436 5228 27488 5234
rect 27172 5166 27200 5199
rect 27436 5170 27488 5176
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27252 5092 27304 5098
rect 27448 5080 27476 5170
rect 27540 5166 27568 6734
rect 29090 6695 29146 6704
rect 28632 6520 28684 6526
rect 28446 6488 28502 6497
rect 28632 6462 28684 6468
rect 28446 6423 28502 6432
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 27620 5296 27672 5302
rect 27620 5238 27672 5244
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27304 5052 27476 5080
rect 27252 5034 27304 5040
rect 27632 4706 27660 5238
rect 27816 5234 27844 5306
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27816 5001 27844 5170
rect 28092 5137 28120 5238
rect 28460 5166 28488 6423
rect 28448 5160 28500 5166
rect 28078 5128 28134 5137
rect 28448 5102 28500 5108
rect 28078 5063 28134 5072
rect 28264 5092 28316 5098
rect 28264 5034 28316 5040
rect 27802 4992 27858 5001
rect 27802 4927 27858 4936
rect 27632 4678 27752 4706
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27632 4146 27660 4558
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27632 3942 27660 4082
rect 27724 3942 27752 4678
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27816 3590 28212 3618
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 27724 3194 27752 3402
rect 27816 3398 27844 3590
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 28000 3398 28028 3470
rect 28184 3466 28212 3590
rect 28172 3460 28224 3466
rect 28172 3402 28224 3408
rect 27804 3392 27856 3398
rect 27804 3334 27856 3340
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27540 2650 27568 2926
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 26976 2100 27028 2106
rect 26976 2042 27028 2048
rect 27448 800 27476 2382
rect 27908 1222 27936 3334
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27988 1420 28040 1426
rect 27988 1362 28040 1368
rect 27896 1216 27948 1222
rect 27896 1158 27948 1164
rect 28000 800 28028 1362
rect 28092 1358 28120 2790
rect 28276 2446 28304 5034
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 28552 3058 28580 4966
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28644 2972 28672 6462
rect 29104 5166 29132 6695
rect 29734 6624 29790 6633
rect 29734 6559 29790 6568
rect 29552 6452 29604 6458
rect 29552 6394 29604 6400
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 28736 3534 28764 4966
rect 29276 4548 29328 4554
rect 29276 4490 29328 4496
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28828 3482 28856 3538
rect 28828 3466 29040 3482
rect 28828 3460 29052 3466
rect 28828 3454 29000 3460
rect 29000 3402 29052 3408
rect 28906 3088 28962 3097
rect 28906 3023 28908 3032
rect 28960 3023 28962 3032
rect 29092 3052 29144 3058
rect 28908 2994 28960 3000
rect 29092 2994 29144 3000
rect 28724 2984 28776 2990
rect 28644 2944 28724 2972
rect 28724 2926 28776 2932
rect 29104 2650 29132 2994
rect 29288 2774 29316 4490
rect 29380 3126 29408 4966
rect 29368 3120 29420 3126
rect 29368 3062 29420 3068
rect 29472 2922 29500 4966
rect 29564 3194 29592 6394
rect 29748 5166 29776 6559
rect 30300 5234 30328 7511
rect 30852 5234 30880 7647
rect 48228 7540 48280 7546
rect 48228 7482 48280 7488
rect 41050 6896 41106 6905
rect 41050 6831 41106 6840
rect 32312 6384 32364 6390
rect 32312 6326 32364 6332
rect 31668 5568 31720 5574
rect 31668 5510 31720 5516
rect 31208 5296 31260 5302
rect 31208 5238 31260 5244
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 29736 5160 29788 5166
rect 29736 5102 29788 5108
rect 30472 5024 30524 5030
rect 29734 4992 29790 5001
rect 30472 4966 30524 4972
rect 29734 4927 29790 4936
rect 29748 4554 29776 4927
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29736 4548 29788 4554
rect 29736 4490 29788 4496
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29656 3058 29684 4422
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29748 3738 29776 4014
rect 29736 3732 29788 3738
rect 29736 3674 29788 3680
rect 30024 3058 30052 4762
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 29460 2916 29512 2922
rect 29460 2858 29512 2864
rect 29288 2746 29500 2774
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28460 1902 28488 2450
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 28540 2304 28592 2310
rect 28540 2246 28592 2252
rect 28552 2038 28580 2246
rect 28540 2032 28592 2038
rect 28540 1974 28592 1980
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 28644 1562 28672 2382
rect 29092 2304 29144 2310
rect 29092 2246 29144 2252
rect 29104 1970 29132 2246
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 28816 1896 28868 1902
rect 28868 1844 29040 1850
rect 28816 1838 29040 1844
rect 28828 1822 29040 1838
rect 29012 1766 29040 1822
rect 29000 1760 29052 1766
rect 29000 1702 29052 1708
rect 28632 1556 28684 1562
rect 28632 1498 28684 1504
rect 28446 1456 28502 1465
rect 28446 1391 28448 1400
rect 28500 1391 28502 1400
rect 28448 1362 28500 1368
rect 28080 1352 28132 1358
rect 29196 1306 29224 2382
rect 29472 1358 29500 2746
rect 29564 1970 29592 2994
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29920 1964 29972 1970
rect 29920 1906 29972 1912
rect 28080 1294 28132 1300
rect 28540 1284 28592 1290
rect 28540 1226 28592 1232
rect 29104 1278 29224 1306
rect 29460 1352 29512 1358
rect 29460 1294 29512 1300
rect 28552 800 28580 1226
rect 29104 800 29132 1278
rect 29656 870 29776 898
rect 29656 800 29684 870
rect 3146 0 3202 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 29748 762 29776 870
rect 29932 762 29960 1906
rect 30208 800 30236 2926
rect 30484 2582 30512 4966
rect 31024 4820 31076 4826
rect 31024 4762 31076 4768
rect 31036 3398 31064 4762
rect 31220 3534 31248 5238
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31404 4690 31432 5170
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31312 4049 31340 4082
rect 31298 4040 31354 4049
rect 31298 3975 31354 3984
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 30932 2984 30984 2990
rect 30932 2926 30984 2932
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30944 2514 30972 2926
rect 31312 2774 31340 3674
rect 31404 3602 31432 4082
rect 31392 3596 31444 3602
rect 31392 3538 31444 3544
rect 31680 3534 31708 5510
rect 31836 4922 32188 5972
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 31836 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 32188 4922
rect 31836 3834 32188 4870
rect 31836 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 32188 3834
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31312 2746 31432 2774
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30300 1902 30328 2246
rect 30288 1896 30340 1902
rect 30288 1838 30340 1844
rect 31036 1562 31064 2382
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31312 1970 31340 2246
rect 31300 1964 31352 1970
rect 31300 1906 31352 1912
rect 31114 1592 31170 1601
rect 31024 1556 31076 1562
rect 31114 1527 31170 1536
rect 31024 1498 31076 1504
rect 31128 1494 31156 1527
rect 31116 1488 31168 1494
rect 31116 1430 31168 1436
rect 30380 1352 30432 1358
rect 30380 1294 30432 1300
rect 29748 734 29960 762
rect 30194 0 30250 800
rect 30392 762 30420 1294
rect 31300 1284 31352 1290
rect 31300 1226 31352 1232
rect 30668 870 30788 898
rect 30668 762 30696 870
rect 30760 800 30788 870
rect 31312 800 31340 1226
rect 31404 1018 31432 2746
rect 31588 2650 31616 2994
rect 31836 2746 32188 3782
rect 32232 3534 32260 5714
rect 32324 3534 32352 6326
rect 34888 6316 34940 6322
rect 34888 6258 34940 6264
rect 33324 5908 33376 5914
rect 33324 5850 33376 5856
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32416 3602 32444 3674
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32218 3088 32274 3097
rect 32600 3058 32628 5714
rect 33048 5024 33100 5030
rect 33048 4966 33100 4972
rect 33060 4214 33088 4966
rect 33048 4208 33100 4214
rect 33048 4150 33100 4156
rect 33048 3528 33100 3534
rect 32692 3476 33048 3482
rect 32692 3470 33100 3476
rect 32692 3454 33088 3470
rect 32692 3398 32720 3454
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 33232 3120 33284 3126
rect 33232 3062 33284 3068
rect 32218 3023 32274 3032
rect 32312 3052 32364 3058
rect 32232 2990 32260 3023
rect 32312 2994 32364 3000
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 33140 3052 33192 3058
rect 33140 2994 33192 3000
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 31836 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 32188 2746
rect 31576 2644 31628 2650
rect 31576 2586 31628 2592
rect 31836 2236 32188 2694
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 31836 2180 31864 2236
rect 31920 2180 31944 2236
rect 32000 2180 32024 2236
rect 32080 2180 32104 2236
rect 32160 2180 32188 2236
rect 31836 2156 32188 2180
rect 31836 2100 31864 2156
rect 31920 2100 31944 2156
rect 32000 2100 32024 2156
rect 32080 2100 32104 2156
rect 32160 2100 32188 2156
rect 31836 2076 32188 2100
rect 31836 2020 31864 2076
rect 31920 2020 31944 2076
rect 32000 2020 32024 2076
rect 32080 2020 32104 2076
rect 32160 2020 32188 2076
rect 31836 1996 32188 2020
rect 31836 1940 31864 1996
rect 31920 1940 31944 1996
rect 32000 1940 32024 1996
rect 32080 1940 32104 1996
rect 32160 1940 32188 1996
rect 31836 1658 32188 1940
rect 31836 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 32188 1658
rect 31836 1040 32188 1606
rect 31392 1012 31444 1018
rect 31392 954 31444 960
rect 31864 870 31984 898
rect 31864 800 31892 870
rect 30392 734 30696 762
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 31956 762 31984 870
rect 32232 762 32260 2382
rect 32324 2106 32352 2994
rect 33152 2650 33180 2994
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 2106 32536 2382
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 32496 2100 32548 2106
rect 32496 2042 32548 2048
rect 32404 1896 32456 1902
rect 32404 1838 32456 1844
rect 32416 800 32444 1838
rect 33244 1358 33272 3062
rect 33336 3058 33364 5850
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33796 4486 33824 4558
rect 33784 4480 33836 4486
rect 33784 4422 33836 4428
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 33428 3194 33456 3674
rect 33416 3188 33468 3194
rect 33416 3130 33468 3136
rect 33796 3058 33824 4082
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 33888 2854 33916 5850
rect 34188 5466 34540 5972
rect 34188 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34540 5466
rect 34058 4856 34114 4865
rect 34058 4791 34114 4800
rect 34072 4622 34100 4791
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 34188 4588 34540 5414
rect 33980 3942 34008 4558
rect 34188 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34540 4588
rect 34188 4508 34540 4532
rect 34188 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34540 4508
rect 34704 4548 34756 4554
rect 34704 4490 34756 4496
rect 34188 4428 34540 4452
rect 34188 4378 34216 4428
rect 34272 4378 34296 4428
rect 34352 4378 34376 4428
rect 34432 4378 34456 4428
rect 34512 4378 34540 4428
rect 34188 4326 34210 4378
rect 34272 4372 34274 4378
rect 34454 4372 34456 4378
rect 34262 4348 34274 4372
rect 34326 4348 34338 4372
rect 34390 4348 34402 4372
rect 34454 4348 34466 4372
rect 34272 4326 34274 4348
rect 34454 4326 34456 4348
rect 34518 4326 34540 4378
rect 34188 4292 34216 4326
rect 34272 4292 34296 4326
rect 34352 4292 34376 4326
rect 34432 4292 34456 4326
rect 34512 4292 34540 4326
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 34188 3290 34540 4292
rect 34716 4146 34744 4490
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 34808 4146 34836 4422
rect 34704 4140 34756 4146
rect 34704 4082 34756 4088
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 34188 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34540 3290
rect 34060 3052 34112 3058
rect 34060 2994 34112 3000
rect 33876 2848 33928 2854
rect 33876 2790 33928 2796
rect 34072 2650 34100 2994
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 32864 1352 32916 1358
rect 32864 1294 32916 1300
rect 33232 1352 33284 1358
rect 33232 1294 33284 1300
rect 32876 950 32904 1294
rect 33048 1284 33100 1290
rect 32968 1244 33048 1272
rect 32864 944 32916 950
rect 32864 886 32916 892
rect 32968 800 32996 1244
rect 33048 1226 33100 1232
rect 33612 1222 33640 2382
rect 34188 2202 34540 3238
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 34188 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34540 2202
rect 34060 1964 34112 1970
rect 34060 1906 34112 1912
rect 33600 1216 33652 1222
rect 33600 1158 33652 1164
rect 33508 944 33560 950
rect 33508 886 33560 892
rect 33520 800 33548 886
rect 34072 800 34100 1906
rect 34188 1114 34540 2150
rect 34624 2106 34652 2994
rect 34612 2100 34664 2106
rect 34612 2042 34664 2048
rect 34704 2100 34756 2106
rect 34704 2042 34756 2048
rect 34612 1896 34664 1902
rect 34612 1838 34664 1844
rect 34188 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34540 1114
rect 34188 1040 34540 1062
rect 34624 800 34652 1838
rect 34716 1766 34744 2042
rect 34808 1970 34836 3062
rect 34900 3058 34928 6258
rect 40406 5808 40462 5817
rect 40406 5743 40462 5752
rect 40420 5710 40448 5743
rect 40408 5704 40460 5710
rect 37002 5672 37058 5681
rect 40408 5646 40460 5652
rect 37002 5607 37004 5616
rect 37056 5607 37058 5616
rect 37004 5578 37056 5584
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35072 4752 35124 4758
rect 35072 4694 35124 4700
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34796 1964 34848 1970
rect 34796 1906 34848 1912
rect 34704 1760 34756 1766
rect 34704 1702 34756 1708
rect 35084 1426 35112 4694
rect 35716 4480 35768 4486
rect 35716 4422 35768 4428
rect 35728 3058 35756 4422
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 35728 2922 35756 2994
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 35912 1834 35940 5510
rect 41064 5370 41092 6831
rect 46388 6520 46440 6526
rect 46388 6462 46440 6468
rect 45652 6248 45704 6254
rect 45652 6190 45704 6196
rect 44916 6180 44968 6186
rect 44916 6122 44968 6128
rect 44638 6080 44694 6089
rect 44638 6015 44694 6024
rect 41512 5704 41564 5710
rect 41512 5646 41564 5652
rect 41694 5672 41750 5681
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 41052 5364 41104 5370
rect 41052 5306 41104 5312
rect 41144 5364 41196 5370
rect 41144 5306 41196 5312
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 3126 36032 3878
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 36832 3058 36860 5306
rect 41156 5250 41184 5306
rect 40972 5234 41184 5250
rect 40960 5228 41184 5234
rect 41012 5222 41184 5228
rect 40960 5170 41012 5176
rect 40408 5160 40460 5166
rect 40408 5102 40460 5108
rect 40420 4010 40448 5102
rect 40592 5092 40644 5098
rect 40592 5034 40644 5040
rect 40604 4826 40632 5034
rect 40592 4820 40644 4826
rect 40592 4762 40644 4768
rect 41236 4616 41288 4622
rect 41236 4558 41288 4564
rect 40408 4004 40460 4010
rect 40408 3946 40460 3952
rect 41248 3670 41276 4558
rect 41236 3664 41288 3670
rect 41236 3606 41288 3612
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 38016 3528 38068 3534
rect 38016 3470 38068 3476
rect 36912 3392 36964 3398
rect 36912 3334 36964 3340
rect 37004 3392 37056 3398
rect 37004 3334 37056 3340
rect 36924 3058 36952 3334
rect 37016 3194 37044 3334
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 36188 2106 36216 2586
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36176 2100 36228 2106
rect 36176 2042 36228 2048
rect 36176 1896 36228 1902
rect 36176 1838 36228 1844
rect 35900 1828 35952 1834
rect 35900 1770 35952 1776
rect 35992 1828 36044 1834
rect 35992 1770 36044 1776
rect 36004 1601 36032 1770
rect 35990 1592 36046 1601
rect 35990 1527 36046 1536
rect 35164 1488 35216 1494
rect 35164 1430 35216 1436
rect 35072 1420 35124 1426
rect 35072 1362 35124 1368
rect 35176 800 35204 1430
rect 35624 1352 35676 1358
rect 35624 1294 35676 1300
rect 35636 1018 35664 1294
rect 36188 1290 36216 1838
rect 36556 1494 36584 2382
rect 36740 2106 36768 2994
rect 36728 2100 36780 2106
rect 36728 2042 36780 2048
rect 37556 1896 37608 1902
rect 37556 1838 37608 1844
rect 37568 1562 37596 1838
rect 37556 1556 37608 1562
rect 37556 1498 37608 1504
rect 36544 1488 36596 1494
rect 36544 1430 36596 1436
rect 37924 1420 37976 1426
rect 37924 1362 37976 1368
rect 37372 1352 37424 1358
rect 37372 1294 37424 1300
rect 36176 1284 36228 1290
rect 36176 1226 36228 1232
rect 36268 1284 36320 1290
rect 36268 1226 36320 1232
rect 35716 1216 35768 1222
rect 35716 1158 35768 1164
rect 35624 1012 35676 1018
rect 35624 954 35676 960
rect 35728 800 35756 1158
rect 36280 800 36308 1226
rect 37384 800 37412 1294
rect 37936 800 37964 1362
rect 38028 1358 38056 3470
rect 39304 2576 39356 2582
rect 39304 2518 39356 2524
rect 39120 2372 39172 2378
rect 39120 2314 39172 2320
rect 39132 2106 39160 2314
rect 39316 2106 39344 2518
rect 39120 2100 39172 2106
rect 39120 2042 39172 2048
rect 39304 2100 39356 2106
rect 39304 2042 39356 2048
rect 39028 1964 39080 1970
rect 39028 1906 39080 1912
rect 38568 1760 38620 1766
rect 38568 1702 38620 1708
rect 38580 1494 38608 1702
rect 38568 1488 38620 1494
rect 38568 1430 38620 1436
rect 38016 1352 38068 1358
rect 38016 1294 38068 1300
rect 39040 800 39068 1906
rect 39776 1358 39804 3538
rect 41418 3360 41474 3369
rect 41418 3295 41474 3304
rect 41432 2446 41460 3295
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41144 1896 41196 1902
rect 41144 1838 41196 1844
rect 41156 1562 41184 1838
rect 41524 1834 41552 5646
rect 41694 5607 41750 5616
rect 41708 5574 41736 5607
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41696 5228 41748 5234
rect 41696 5170 41748 5176
rect 41708 4758 41736 5170
rect 41836 4922 42188 5972
rect 43812 5704 43864 5710
rect 43812 5646 43864 5652
rect 42708 5160 42760 5166
rect 42706 5128 42708 5137
rect 42760 5128 42762 5137
rect 42706 5063 42762 5072
rect 41836 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 42188 4922
rect 41696 4752 41748 4758
rect 41696 4694 41748 4700
rect 41696 4616 41748 4622
rect 41696 4558 41748 4564
rect 41708 4078 41736 4558
rect 41696 4072 41748 4078
rect 41696 4014 41748 4020
rect 41836 3834 42188 4870
rect 43352 4684 43404 4690
rect 43352 4626 43404 4632
rect 42524 4480 42576 4486
rect 42524 4422 42576 4428
rect 42616 4480 42668 4486
rect 42616 4422 42668 4428
rect 42536 4010 42564 4422
rect 42628 4078 42656 4422
rect 43364 4185 43392 4626
rect 43536 4616 43588 4622
rect 43536 4558 43588 4564
rect 43350 4176 43406 4185
rect 43350 4111 43406 4120
rect 42616 4072 42668 4078
rect 42616 4014 42668 4020
rect 42524 4004 42576 4010
rect 42524 3946 42576 3952
rect 41836 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 42188 3834
rect 41836 2746 42188 3782
rect 42248 3664 42300 3670
rect 42248 3606 42300 3612
rect 41836 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 42188 2746
rect 41836 2236 42188 2694
rect 41836 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 42188 2236
rect 41836 2156 42188 2180
rect 41696 2100 41748 2106
rect 41696 2042 41748 2048
rect 41836 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 42188 2156
rect 42260 2106 42288 3606
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42340 2440 42392 2446
rect 42340 2382 42392 2388
rect 41836 2076 42188 2100
rect 41512 1828 41564 1834
rect 41512 1770 41564 1776
rect 41144 1556 41196 1562
rect 41144 1498 41196 1504
rect 41708 1494 41736 2042
rect 41836 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 42188 2076
rect 42248 2100 42300 2106
rect 42248 2042 42300 2048
rect 41836 1996 42188 2020
rect 41836 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 42188 1996
rect 41836 1658 42188 1940
rect 41836 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 42188 1658
rect 41696 1488 41748 1494
rect 41696 1430 41748 1436
rect 41236 1420 41288 1426
rect 41236 1362 41288 1368
rect 39764 1352 39816 1358
rect 40776 1352 40828 1358
rect 39764 1294 39816 1300
rect 40696 1312 40776 1340
rect 39580 1284 39632 1290
rect 39580 1226 39632 1232
rect 39592 800 39620 1226
rect 40696 800 40724 1312
rect 40776 1294 40828 1300
rect 41248 800 41276 1362
rect 41836 1040 42188 1606
rect 42352 800 42380 2382
rect 42444 1358 42472 2994
rect 42984 2984 43036 2990
rect 42984 2926 43036 2932
rect 42996 1970 43024 2926
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 42892 1964 42944 1970
rect 42892 1906 42944 1912
rect 42984 1964 43036 1970
rect 42984 1906 43036 1912
rect 42904 1358 42932 1906
rect 42984 1828 43036 1834
rect 42984 1770 43036 1776
rect 42432 1352 42484 1358
rect 42432 1294 42484 1300
rect 42892 1352 42944 1358
rect 42892 1294 42944 1300
rect 42996 1034 43024 1770
rect 42904 1006 43024 1034
rect 42904 800 42932 1006
rect 43456 800 43484 2382
rect 43548 2310 43576 4558
rect 43536 2304 43588 2310
rect 43536 2246 43588 2252
rect 43824 882 43852 5646
rect 44188 5466 44540 5972
rect 44652 5710 44680 6015
rect 44928 5710 44956 6122
rect 45664 5710 45692 6190
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46308 5710 46336 6054
rect 46400 5710 46428 6462
rect 47492 6452 47544 6458
rect 47492 6394 47544 6400
rect 46754 6216 46810 6225
rect 46754 6151 46810 6160
rect 47032 6180 47084 6186
rect 44640 5704 44692 5710
rect 44640 5646 44692 5652
rect 44916 5704 44968 5710
rect 44916 5646 44968 5652
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 46296 5704 46348 5710
rect 46296 5646 46348 5652
rect 46388 5704 46440 5710
rect 46388 5646 46440 5652
rect 44188 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 44540 5466
rect 44188 4588 44540 5414
rect 46202 5400 46258 5409
rect 46202 5335 46258 5344
rect 46216 5234 46244 5335
rect 46204 5228 46256 5234
rect 46204 5170 46256 5176
rect 46296 5228 46348 5234
rect 46296 5170 46348 5176
rect 44640 5092 44692 5098
rect 44640 5034 44692 5040
rect 44188 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 44540 4588
rect 44188 4508 44540 4532
rect 43996 4480 44048 4486
rect 43996 4422 44048 4428
rect 44188 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 44540 4508
rect 44188 4428 44540 4452
rect 44008 4214 44036 4422
rect 44188 4378 44216 4428
rect 44272 4378 44296 4428
rect 44352 4378 44376 4428
rect 44432 4378 44456 4428
rect 44512 4378 44540 4428
rect 44188 4326 44210 4378
rect 44272 4372 44274 4378
rect 44454 4372 44456 4378
rect 44262 4348 44274 4372
rect 44326 4348 44338 4372
rect 44390 4348 44402 4372
rect 44454 4348 44466 4372
rect 44272 4326 44274 4348
rect 44454 4326 44456 4348
rect 44518 4326 44540 4378
rect 44188 4292 44216 4326
rect 44272 4292 44296 4326
rect 44352 4292 44376 4326
rect 44432 4292 44456 4326
rect 44512 4292 44540 4326
rect 43996 4208 44048 4214
rect 43996 4150 44048 4156
rect 44188 3290 44540 4292
rect 44652 3466 44680 5034
rect 46020 5024 46072 5030
rect 44730 4992 44786 5001
rect 46020 4966 46072 4972
rect 44730 4927 44786 4936
rect 44744 4826 44772 4927
rect 46032 4826 46060 4966
rect 44732 4820 44784 4826
rect 44732 4762 44784 4768
rect 46020 4820 46072 4826
rect 46020 4762 46072 4768
rect 45100 4752 45152 4758
rect 45100 4694 45152 4700
rect 44732 4684 44784 4690
rect 44732 4626 44784 4632
rect 44744 4185 44772 4626
rect 44730 4176 44786 4185
rect 44730 4111 44786 4120
rect 45112 4010 45140 4694
rect 46308 4622 46336 5170
rect 46572 5160 46624 5166
rect 46572 5102 46624 5108
rect 46296 4616 46348 4622
rect 46296 4558 46348 4564
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 45100 4004 45152 4010
rect 45100 3946 45152 3952
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 44640 3460 44692 3466
rect 44640 3402 44692 3408
rect 44188 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 44540 3290
rect 44188 2202 44540 3238
rect 44836 2922 44864 3470
rect 45940 3058 45968 4422
rect 45928 3052 45980 3058
rect 45928 2994 45980 3000
rect 44824 2916 44876 2922
rect 44824 2858 44876 2864
rect 44732 2576 44784 2582
rect 44732 2518 44784 2524
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44188 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 44540 2202
rect 43996 1284 44048 1290
rect 43996 1226 44048 1232
rect 43812 876 43864 882
rect 43812 818 43864 824
rect 44008 800 44036 1226
rect 44188 1114 44540 2150
rect 44652 1426 44680 2314
rect 44640 1420 44692 1426
rect 44640 1362 44692 1368
rect 44744 1358 44772 2518
rect 44836 2106 44864 2858
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44824 2100 44876 2106
rect 44824 2042 44876 2048
rect 44824 1420 44876 1426
rect 44824 1362 44876 1368
rect 44732 1352 44784 1358
rect 44732 1294 44784 1300
rect 44188 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 44540 1114
rect 44188 1040 44540 1062
rect 44560 870 44680 898
rect 44560 800 44588 870
rect 31956 734 32260 762
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 44652 762 44680 870
rect 44836 762 44864 1362
rect 44928 1358 44956 2790
rect 46584 2650 46612 5102
rect 46768 4622 46796 6151
rect 47032 6122 47084 6128
rect 47044 5710 47072 6122
rect 47504 5710 47532 6394
rect 48136 6384 48188 6390
rect 48136 6326 48188 6332
rect 47032 5704 47084 5710
rect 47032 5646 47084 5652
rect 47492 5704 47544 5710
rect 47492 5646 47544 5652
rect 47872 5642 48084 5658
rect 47860 5636 48096 5642
rect 47912 5630 48044 5636
rect 47860 5578 47912 5584
rect 48044 5578 48096 5584
rect 48148 5574 48176 6326
rect 48136 5568 48188 5574
rect 48136 5510 48188 5516
rect 48240 5166 48268 7482
rect 48872 6860 48924 6866
rect 48872 6802 48924 6808
rect 48884 5778 48912 6802
rect 49608 6452 49660 6458
rect 49608 6394 49660 6400
rect 49620 5914 49648 6394
rect 51080 6248 51132 6254
rect 51080 6190 51132 6196
rect 48964 5908 49016 5914
rect 48964 5850 49016 5856
rect 49608 5908 49660 5914
rect 49608 5850 49660 5856
rect 48976 5778 49004 5850
rect 48872 5772 48924 5778
rect 48872 5714 48924 5720
rect 48964 5772 49016 5778
rect 48964 5714 49016 5720
rect 50436 5704 50488 5710
rect 50436 5646 50488 5652
rect 48962 5536 49018 5545
rect 48962 5471 49018 5480
rect 47492 5160 47544 5166
rect 47228 5098 47440 5114
rect 47492 5102 47544 5108
rect 48228 5160 48280 5166
rect 48228 5102 48280 5108
rect 47216 5092 47452 5098
rect 47268 5086 47400 5092
rect 47216 5034 47268 5040
rect 47400 5034 47452 5040
rect 47124 5024 47176 5030
rect 47124 4966 47176 4972
rect 46664 4616 46716 4622
rect 46664 4558 46716 4564
rect 46756 4616 46808 4622
rect 46756 4558 46808 4564
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46676 4468 46704 4558
rect 46860 4468 46888 4558
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 46676 4440 46888 4468
rect 46952 4078 46980 4490
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 47032 3120 47084 3126
rect 47032 3062 47084 3068
rect 46572 2644 46624 2650
rect 46572 2586 46624 2592
rect 45560 2440 45612 2446
rect 45560 2382 45612 2388
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 45468 2100 45520 2106
rect 45468 2042 45520 2048
rect 45480 1562 45508 2042
rect 45572 1562 45600 2382
rect 45652 1964 45704 1970
rect 45652 1906 45704 1912
rect 45468 1556 45520 1562
rect 45468 1498 45520 1504
rect 45560 1556 45612 1562
rect 45560 1498 45612 1504
rect 44916 1352 44968 1358
rect 44916 1294 44968 1300
rect 45100 1284 45152 1290
rect 45100 1226 45152 1232
rect 45112 800 45140 1226
rect 45664 800 45692 1906
rect 46216 1902 46244 2382
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 46860 1970 46888 2246
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46020 1896 46072 1902
rect 46020 1838 46072 1844
rect 46204 1896 46256 1902
rect 46204 1838 46256 1844
rect 46032 1222 46060 1838
rect 46940 1828 46992 1834
rect 46940 1770 46992 1776
rect 46952 1562 46980 1770
rect 46940 1556 46992 1562
rect 46940 1498 46992 1504
rect 47044 1494 47072 3062
rect 47136 3058 47164 4966
rect 47504 3738 47532 5102
rect 48976 4690 49004 5471
rect 49148 5160 49200 5166
rect 49148 5102 49200 5108
rect 48964 4684 49016 4690
rect 48964 4626 49016 4632
rect 49056 4480 49108 4486
rect 49056 4422 49108 4428
rect 47492 3732 47544 3738
rect 47492 3674 47544 3680
rect 48228 3460 48280 3466
rect 48228 3402 48280 3408
rect 47492 3392 47544 3398
rect 47492 3334 47544 3340
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 47216 2576 47268 2582
rect 47216 2518 47268 2524
rect 47228 1766 47256 2518
rect 47308 2440 47360 2446
rect 47308 2382 47360 2388
rect 47216 1760 47268 1766
rect 47216 1702 47268 1708
rect 47032 1488 47084 1494
rect 47032 1430 47084 1436
rect 46204 1420 46256 1426
rect 46204 1362 46256 1368
rect 46020 1216 46072 1222
rect 46020 1158 46072 1164
rect 46216 800 46244 1362
rect 47320 800 47348 2382
rect 47504 1358 47532 3334
rect 47584 2848 47636 2854
rect 47584 2790 47636 2796
rect 47596 1970 47624 2790
rect 48240 2650 48268 3402
rect 49068 3058 49096 4422
rect 49160 3942 49188 5102
rect 49516 5024 49568 5030
rect 49516 4966 49568 4972
rect 49424 4616 49476 4622
rect 49424 4558 49476 4564
rect 49436 4214 49464 4558
rect 49528 4214 49556 4966
rect 49424 4208 49476 4214
rect 49424 4150 49476 4156
rect 49516 4208 49568 4214
rect 49516 4150 49568 4156
rect 49148 3936 49200 3942
rect 49148 3878 49200 3884
rect 49056 3052 49108 3058
rect 49056 2994 49108 3000
rect 50068 2916 50120 2922
rect 50068 2858 50120 2864
rect 48228 2644 48280 2650
rect 48228 2586 48280 2592
rect 48872 2440 48924 2446
rect 48872 2382 48924 2388
rect 48964 2440 49016 2446
rect 48964 2382 49016 2388
rect 47584 1964 47636 1970
rect 47584 1906 47636 1912
rect 47860 1896 47912 1902
rect 47860 1838 47912 1844
rect 47492 1352 47544 1358
rect 47492 1294 47544 1300
rect 47872 800 47900 1838
rect 48884 1358 48912 2382
rect 48872 1352 48924 1358
rect 48872 1294 48924 1300
rect 48976 800 49004 2382
rect 49424 2304 49476 2310
rect 49424 2246 49476 2252
rect 49516 2304 49568 2310
rect 49516 2246 49568 2252
rect 49436 1358 49464 2246
rect 49528 1970 49556 2246
rect 49516 1964 49568 1970
rect 49516 1906 49568 1912
rect 49608 1420 49660 1426
rect 49528 1380 49608 1408
rect 49424 1352 49476 1358
rect 49424 1294 49476 1300
rect 49528 800 49556 1380
rect 49608 1362 49660 1368
rect 50080 1358 50108 2858
rect 50448 2106 50476 5646
rect 51092 5522 51120 6190
rect 51264 5704 51316 5710
rect 51264 5646 51316 5652
rect 51000 5494 51120 5522
rect 51000 5166 51028 5494
rect 50988 5160 51040 5166
rect 50988 5102 51040 5108
rect 51276 3126 51304 5646
rect 51836 4922 52188 5972
rect 52288 5710 52316 7686
rect 56140 7676 56192 7682
rect 56140 7618 56192 7624
rect 55588 6996 55640 7002
rect 55588 6938 55640 6944
rect 54668 6520 54720 6526
rect 54668 6462 54720 6468
rect 53932 6316 53984 6322
rect 53932 6258 53984 6264
rect 53944 5710 53972 6258
rect 52276 5704 52328 5710
rect 52276 5646 52328 5652
rect 52644 5704 52696 5710
rect 52644 5646 52696 5652
rect 53380 5704 53432 5710
rect 53380 5646 53432 5652
rect 53932 5704 53984 5710
rect 53932 5646 53984 5652
rect 51836 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 52188 4922
rect 51836 3834 52188 4870
rect 51836 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 52188 3834
rect 51540 3596 51592 3602
rect 51540 3538 51592 3544
rect 51264 3120 51316 3126
rect 51264 3062 51316 3068
rect 51552 2106 51580 3538
rect 51836 2746 52188 3782
rect 52656 3670 52684 5646
rect 53012 5228 53064 5234
rect 53012 5170 53064 5176
rect 52920 5024 52972 5030
rect 52920 4966 52972 4972
rect 52644 3664 52696 3670
rect 52644 3606 52696 3612
rect 52932 3058 52960 4966
rect 53024 4758 53052 5170
rect 53288 5160 53340 5166
rect 53288 5102 53340 5108
rect 53012 4752 53064 4758
rect 53012 4694 53064 4700
rect 53300 4214 53328 5102
rect 53288 4208 53340 4214
rect 53288 4150 53340 4156
rect 52920 3052 52972 3058
rect 52920 2994 52972 3000
rect 52644 2848 52696 2854
rect 52644 2790 52696 2796
rect 53104 2848 53156 2854
rect 53104 2790 53156 2796
rect 51836 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 52188 2746
rect 51836 2236 52188 2694
rect 51836 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 52188 2236
rect 51836 2156 52188 2180
rect 50436 2100 50488 2106
rect 50436 2042 50488 2048
rect 51540 2100 51592 2106
rect 51540 2042 51592 2048
rect 51836 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 52188 2156
rect 51836 2076 52188 2100
rect 51836 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 52188 2076
rect 51836 1996 52188 2020
rect 51836 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 52188 1996
rect 51264 1896 51316 1902
rect 51264 1838 51316 1844
rect 51276 1562 51304 1838
rect 51836 1658 52188 1940
rect 51836 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 52188 1658
rect 51264 1556 51316 1562
rect 51264 1498 51316 1504
rect 50068 1352 50120 1358
rect 50068 1294 50120 1300
rect 50620 1352 50672 1358
rect 50620 1294 50672 1300
rect 50632 800 50660 1294
rect 51172 1284 51224 1290
rect 51172 1226 51224 1232
rect 51184 800 51212 1226
rect 51836 1040 52188 1606
rect 52656 1358 52684 2790
rect 53116 1970 53144 2790
rect 53104 1964 53156 1970
rect 53104 1906 53156 1912
rect 52828 1896 52880 1902
rect 52828 1838 52880 1844
rect 52644 1352 52696 1358
rect 52644 1294 52696 1300
rect 52276 1216 52328 1222
rect 52276 1158 52328 1164
rect 52288 800 52316 1158
rect 52840 800 52868 1838
rect 53392 1766 53420 5646
rect 54188 5466 54540 5944
rect 54680 5778 54708 6462
rect 55600 6254 55628 6938
rect 55680 6928 55732 6934
rect 55680 6870 55732 6876
rect 55588 6248 55640 6254
rect 55588 6190 55640 6196
rect 55692 5914 55720 6870
rect 56048 6860 56100 6866
rect 56048 6802 56100 6808
rect 55862 6352 55918 6361
rect 55862 6287 55918 6296
rect 55772 6180 55824 6186
rect 55772 6122 55824 6128
rect 55784 5914 55812 6122
rect 55876 6089 55904 6287
rect 56060 6186 56088 6802
rect 56048 6180 56100 6186
rect 56048 6122 56100 6128
rect 55956 6112 56008 6118
rect 55862 6080 55918 6089
rect 55956 6054 56008 6060
rect 55862 6015 55918 6024
rect 55680 5908 55732 5914
rect 55680 5850 55732 5856
rect 55772 5908 55824 5914
rect 55772 5850 55824 5856
rect 55968 5846 55996 6054
rect 55956 5840 56008 5846
rect 55956 5782 56008 5788
rect 54668 5772 54720 5778
rect 54668 5714 54720 5720
rect 56152 5710 56180 7618
rect 56508 7608 56560 7614
rect 56508 7550 56560 7556
rect 56232 5840 56284 5846
rect 56232 5782 56284 5788
rect 54576 5704 54628 5710
rect 54576 5646 54628 5652
rect 55312 5704 55364 5710
rect 55312 5646 55364 5652
rect 56140 5704 56192 5710
rect 56140 5646 56192 5652
rect 54188 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 54540 5466
rect 54188 4588 54540 5414
rect 54188 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 54540 4588
rect 54188 4508 54540 4532
rect 54188 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 54540 4508
rect 54188 4428 54540 4452
rect 54188 4378 54216 4428
rect 54272 4378 54296 4428
rect 54352 4378 54376 4428
rect 54432 4378 54456 4428
rect 54512 4378 54540 4428
rect 54188 4326 54210 4378
rect 54272 4372 54274 4378
rect 54454 4372 54456 4378
rect 54262 4348 54274 4372
rect 54326 4348 54338 4372
rect 54390 4348 54402 4372
rect 54454 4348 54466 4372
rect 54272 4326 54274 4348
rect 54454 4326 54456 4348
rect 54518 4326 54540 4378
rect 54188 4292 54216 4326
rect 54272 4292 54296 4326
rect 54352 4292 54376 4326
rect 54432 4292 54456 4326
rect 54512 4292 54540 4326
rect 54024 4004 54076 4010
rect 54024 3946 54076 3952
rect 53932 3052 53984 3058
rect 53932 2994 53984 3000
rect 53944 2650 53972 2994
rect 53932 2644 53984 2650
rect 53932 2586 53984 2592
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53932 2440 53984 2446
rect 53932 2382 53984 2388
rect 53380 1760 53432 1766
rect 53380 1702 53432 1708
rect 53852 1358 53880 2382
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 53944 800 53972 2382
rect 54036 2378 54064 3946
rect 54188 3290 54540 4292
rect 54588 4010 54616 5646
rect 54680 5494 55076 5522
rect 54680 5302 54708 5494
rect 54760 5364 54812 5370
rect 54760 5306 54812 5312
rect 54668 5296 54720 5302
rect 54668 5238 54720 5244
rect 54772 5148 54800 5306
rect 55048 5302 55076 5494
rect 55036 5296 55088 5302
rect 55036 5238 55088 5244
rect 55128 5160 55180 5166
rect 54772 5120 55128 5148
rect 55128 5102 55180 5108
rect 54668 5024 54720 5030
rect 54668 4966 54720 4972
rect 54576 4004 54628 4010
rect 54576 3946 54628 3952
rect 54188 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 54540 3290
rect 54024 2372 54076 2378
rect 54024 2314 54076 2320
rect 54188 2202 54540 3238
rect 54680 3058 54708 4966
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 55220 2848 55272 2854
rect 55220 2790 55272 2796
rect 55036 2372 55088 2378
rect 55036 2314 55088 2320
rect 54760 2304 54812 2310
rect 54760 2246 54812 2252
rect 54188 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 54540 2202
rect 54188 1114 54540 2150
rect 54772 1970 54800 2246
rect 55048 2106 55076 2314
rect 55036 2100 55088 2106
rect 55036 2042 55088 2048
rect 54760 1964 54812 1970
rect 54760 1906 54812 1912
rect 55232 1358 55260 2790
rect 55324 2582 55352 5646
rect 55954 5536 56010 5545
rect 55954 5471 56010 5480
rect 55968 5098 55996 5471
rect 55956 5092 56008 5098
rect 55956 5034 56008 5040
rect 55772 3664 55824 3670
rect 55772 3606 55824 3612
rect 55312 2576 55364 2582
rect 55312 2518 55364 2524
rect 55588 1896 55640 1902
rect 55588 1838 55640 1844
rect 55220 1352 55272 1358
rect 55220 1294 55272 1300
rect 54576 1284 54628 1290
rect 54576 1226 54628 1232
rect 54188 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 54540 1114
rect 54188 1040 54540 1062
rect 54588 898 54616 1226
rect 54496 870 54616 898
rect 54496 800 54524 870
rect 55600 800 55628 1838
rect 55784 1834 55812 3606
rect 56244 3058 56272 5782
rect 56520 5778 56548 7550
rect 59188 7478 59216 7772
rect 59560 7754 59612 7760
rect 59176 7472 59228 7478
rect 59176 7414 59228 7420
rect 60372 7268 60424 7274
rect 60372 7210 60424 7216
rect 60096 7064 60148 7070
rect 60096 7006 60148 7012
rect 60004 6860 60056 6866
rect 60004 6802 60056 6808
rect 59544 6520 59596 6526
rect 59544 6462 59596 6468
rect 59636 6520 59688 6526
rect 59636 6462 59688 6468
rect 58162 5944 58218 5953
rect 58162 5879 58218 5888
rect 58176 5778 58204 5879
rect 56508 5772 56560 5778
rect 56508 5714 56560 5720
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 58164 5772 58216 5778
rect 58164 5714 58216 5720
rect 58256 5772 58308 5778
rect 58256 5714 58308 5720
rect 56324 5704 56376 5710
rect 56324 5646 56376 5652
rect 56336 5234 56364 5646
rect 56324 5228 56376 5234
rect 56324 5170 56376 5176
rect 56416 5228 56468 5234
rect 56416 5170 56468 5176
rect 56428 4146 56456 5170
rect 56416 4140 56468 4146
rect 56416 4082 56468 4088
rect 57808 3058 57836 5714
rect 58268 5574 58296 5714
rect 59556 5574 59584 6462
rect 59648 5778 59676 6462
rect 60016 6322 60044 6802
rect 59912 6316 59964 6322
rect 59912 6258 59964 6264
rect 60004 6316 60056 6322
rect 60004 6258 60056 6264
rect 59726 6080 59782 6089
rect 59726 6015 59782 6024
rect 59740 5778 59768 6015
rect 59924 5914 59952 6258
rect 59820 5908 59872 5914
rect 59820 5850 59872 5856
rect 59912 5908 59964 5914
rect 59912 5850 59964 5856
rect 59832 5778 59860 5850
rect 59636 5772 59688 5778
rect 59636 5714 59688 5720
rect 59728 5772 59780 5778
rect 59728 5714 59780 5720
rect 59820 5772 59872 5778
rect 59820 5714 59872 5720
rect 58256 5568 58308 5574
rect 58256 5510 58308 5516
rect 59452 5568 59504 5574
rect 59452 5510 59504 5516
rect 59544 5568 59596 5574
rect 59544 5510 59596 5516
rect 58532 3732 58584 3738
rect 58532 3674 58584 3680
rect 58544 3534 58572 3674
rect 58532 3528 58584 3534
rect 58532 3470 58584 3476
rect 59464 3058 59492 5510
rect 60108 4826 60136 7006
rect 60096 4820 60148 4826
rect 60096 4762 60148 4768
rect 60384 4758 60412 7210
rect 61566 7032 61622 7041
rect 61566 6967 61622 6976
rect 61476 5840 61528 5846
rect 61580 5817 61608 6967
rect 61476 5782 61528 5788
rect 61566 5808 61622 5817
rect 61108 5704 61160 5710
rect 61108 5646 61160 5652
rect 61016 5636 61068 5642
rect 61016 5578 61068 5584
rect 61028 5545 61056 5578
rect 61014 5536 61070 5545
rect 61014 5471 61070 5480
rect 60648 5364 60700 5370
rect 60648 5306 60700 5312
rect 60372 4752 60424 4758
rect 60372 4694 60424 4700
rect 60660 4185 60688 5306
rect 61120 4826 61148 5646
rect 61488 5574 61516 5782
rect 61672 5778 61700 7822
rect 62488 7812 62540 7818
rect 62488 7754 62540 7760
rect 62302 6624 62358 6633
rect 62500 6594 62528 7754
rect 63420 7682 63448 10286
rect 63512 7886 63540 67712
rect 63592 60920 63644 60926
rect 63592 60862 63644 60868
rect 63500 7880 63552 7886
rect 63500 7822 63552 7828
rect 63408 7676 63460 7682
rect 63408 7618 63460 7624
rect 63604 7614 63632 60862
rect 63696 17921 63724 69566
rect 64892 68950 64920 71062
rect 64880 68944 64932 68950
rect 64880 68886 64932 68892
rect 64880 66496 64932 66502
rect 64880 66438 64932 66444
rect 64892 64326 64920 66438
rect 64880 64320 64932 64326
rect 64880 64262 64932 64268
rect 64892 62150 64920 64262
rect 64880 62144 64932 62150
rect 64880 62086 64932 62092
rect 64892 60314 64920 62086
rect 64880 60308 64932 60314
rect 64880 60250 64932 60256
rect 64892 58070 64920 60250
rect 64880 58064 64932 58070
rect 64880 58006 64932 58012
rect 64892 55622 64920 58006
rect 64880 55616 64932 55622
rect 64880 55558 64932 55564
rect 64892 53582 64920 55558
rect 64880 53576 64932 53582
rect 64880 53518 64932 53524
rect 63774 52592 63830 52601
rect 63774 52527 63830 52536
rect 63788 52494 63816 52527
rect 63776 52488 63828 52494
rect 63776 52430 63828 52436
rect 64892 51542 64920 53518
rect 64880 51536 64932 51542
rect 64880 51478 64932 51484
rect 63776 50312 63828 50318
rect 63774 50280 63776 50289
rect 63828 50280 63830 50289
rect 63774 50215 63830 50224
rect 64972 48136 65024 48142
rect 64970 48104 64972 48113
rect 65024 48104 65026 48113
rect 64970 48039 65026 48048
rect 64420 47728 64472 47734
rect 64418 47696 64420 47705
rect 64472 47696 64474 47705
rect 64418 47631 64474 47640
rect 64604 47388 64656 47394
rect 64604 47330 64656 47336
rect 63868 47048 63920 47054
rect 63868 46990 63920 46996
rect 63774 43344 63830 43353
rect 63774 43279 63776 43288
rect 63828 43279 63830 43288
rect 63776 43250 63828 43256
rect 63776 25288 63828 25294
rect 63776 25230 63828 25236
rect 63682 17912 63738 17921
rect 63682 17847 63738 17856
rect 63684 16584 63736 16590
rect 63684 16526 63736 16532
rect 63696 11914 63724 16526
rect 63788 12050 63816 25230
rect 63880 12186 63908 46990
rect 64052 45960 64104 45966
rect 64052 45902 64104 45908
rect 63960 45280 64012 45286
rect 63960 45222 64012 45228
rect 63972 12306 64000 45222
rect 63960 12300 64012 12306
rect 63960 12242 64012 12248
rect 63880 12158 64000 12186
rect 63788 12022 63908 12050
rect 63696 11886 63816 11914
rect 63682 11792 63738 11801
rect 63682 11727 63738 11736
rect 63696 7750 63724 11727
rect 63684 7744 63736 7750
rect 63684 7686 63736 7692
rect 63592 7608 63644 7614
rect 63592 7550 63644 7556
rect 62764 7404 62816 7410
rect 62764 7346 62816 7352
rect 62302 6559 62358 6568
rect 62488 6588 62540 6594
rect 62316 6225 62344 6559
rect 62488 6530 62540 6536
rect 61750 6216 61806 6225
rect 61750 6151 61806 6160
rect 62302 6216 62358 6225
rect 62302 6151 62358 6160
rect 61764 5817 61792 6151
rect 61750 5808 61806 5817
rect 61566 5743 61622 5752
rect 61660 5772 61712 5778
rect 61750 5743 61806 5752
rect 61660 5714 61712 5720
rect 61200 5568 61252 5574
rect 61200 5510 61252 5516
rect 61476 5568 61528 5574
rect 61476 5510 61528 5516
rect 61108 4820 61160 4826
rect 61108 4762 61160 4768
rect 60752 4554 60964 4570
rect 60740 4548 60964 4554
rect 60792 4542 60964 4548
rect 60740 4490 60792 4496
rect 60832 4480 60884 4486
rect 60936 4468 60964 4542
rect 61016 4480 61068 4486
rect 60936 4440 61016 4468
rect 60832 4422 60884 4428
rect 61016 4422 61068 4428
rect 60646 4176 60702 4185
rect 60646 4111 60702 4120
rect 60844 4010 60872 4422
rect 61108 4140 61160 4146
rect 61108 4082 61160 4088
rect 60832 4004 60884 4010
rect 60832 3946 60884 3952
rect 60740 3528 60792 3534
rect 60740 3470 60792 3476
rect 56232 3052 56284 3058
rect 56232 2994 56284 3000
rect 57796 3052 57848 3058
rect 57796 2994 57848 3000
rect 59452 3052 59504 3058
rect 59452 2994 59504 3000
rect 56416 2848 56468 2854
rect 56416 2790 56468 2796
rect 57980 2848 58032 2854
rect 57980 2790 58032 2796
rect 60372 2848 60424 2854
rect 60372 2790 60424 2796
rect 56428 1970 56456 2790
rect 57336 2440 57388 2446
rect 57336 2382 57388 2388
rect 56692 2372 56744 2378
rect 56692 2314 56744 2320
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 56140 1896 56192 1902
rect 56140 1838 56192 1844
rect 55772 1828 55824 1834
rect 55772 1770 55824 1776
rect 56152 800 56180 1838
rect 56704 1358 56732 2314
rect 57244 1760 57296 1766
rect 57244 1702 57296 1708
rect 57256 1358 57284 1702
rect 56692 1352 56744 1358
rect 56692 1294 56744 1300
rect 57244 1352 57296 1358
rect 57244 1294 57296 1300
rect 57348 1170 57376 2382
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 57900 1970 57928 2246
rect 57888 1964 57940 1970
rect 57888 1906 57940 1912
rect 57992 1358 58020 2790
rect 59360 1896 59412 1902
rect 59360 1838 59412 1844
rect 59372 1358 59400 1838
rect 59452 1420 59504 1426
rect 59452 1362 59504 1368
rect 57980 1352 58032 1358
rect 57980 1294 58032 1300
rect 59360 1352 59412 1358
rect 59360 1294 59412 1300
rect 57796 1284 57848 1290
rect 57796 1226 57848 1232
rect 58900 1284 58952 1290
rect 58900 1226 58952 1232
rect 57256 1142 57376 1170
rect 57256 800 57284 1142
rect 57808 800 57836 1226
rect 58912 800 58940 1226
rect 59464 800 59492 1362
rect 60384 1358 60412 2790
rect 60752 2650 60780 3470
rect 60740 2644 60792 2650
rect 60740 2586 60792 2592
rect 61016 2372 61068 2378
rect 61016 2314 61068 2320
rect 60556 1896 60608 1902
rect 60556 1838 60608 1844
rect 60372 1352 60424 1358
rect 60372 1294 60424 1300
rect 60568 800 60596 1838
rect 61028 1562 61056 2314
rect 61120 2106 61148 4082
rect 61212 3058 61240 5510
rect 61292 5228 61344 5234
rect 61292 5170 61344 5176
rect 61304 4622 61332 5170
rect 61836 4922 62188 5972
rect 62776 5953 62804 7346
rect 63040 7336 63092 7342
rect 63040 7278 63092 7284
rect 62946 6896 63002 6905
rect 62946 6831 63002 6840
rect 62762 5944 62818 5953
rect 62762 5879 62818 5888
rect 62960 5778 62988 6831
rect 63052 6118 63080 7278
rect 63500 6588 63552 6594
rect 63500 6530 63552 6536
rect 63040 6112 63092 6118
rect 63040 6054 63092 6060
rect 63132 6112 63184 6118
rect 63132 6054 63184 6060
rect 63040 5908 63092 5914
rect 63040 5850 63092 5856
rect 63052 5778 63080 5850
rect 62948 5772 63000 5778
rect 62948 5714 63000 5720
rect 63040 5772 63092 5778
rect 63040 5714 63092 5720
rect 63144 5574 63172 6054
rect 63316 5908 63368 5914
rect 63316 5850 63368 5856
rect 63132 5568 63184 5574
rect 63132 5510 63184 5516
rect 63224 5568 63276 5574
rect 63224 5510 63276 5516
rect 61836 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 62188 4922
rect 61384 4684 61436 4690
rect 61384 4626 61436 4632
rect 61292 4616 61344 4622
rect 61292 4558 61344 4564
rect 61304 3738 61332 4558
rect 61396 4185 61424 4626
rect 61382 4176 61438 4185
rect 61382 4111 61438 4120
rect 61836 3834 62188 4870
rect 62672 4752 62724 4758
rect 62672 4694 62724 4700
rect 62684 4622 62712 4694
rect 62672 4616 62724 4622
rect 62672 4558 62724 4564
rect 62764 4548 62816 4554
rect 62764 4490 62816 4496
rect 62776 4010 62804 4490
rect 62764 4004 62816 4010
rect 62764 3946 62816 3952
rect 61836 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 62188 3834
rect 61292 3732 61344 3738
rect 61292 3674 61344 3680
rect 61200 3052 61252 3058
rect 61200 2994 61252 3000
rect 61384 2848 61436 2854
rect 61384 2790 61436 2796
rect 61108 2100 61160 2106
rect 61108 2042 61160 2048
rect 61396 1970 61424 2790
rect 61836 2746 62188 3782
rect 63236 3058 63264 5510
rect 63328 5273 63356 5850
rect 63408 5568 63460 5574
rect 63406 5536 63408 5545
rect 63460 5536 63462 5545
rect 63406 5471 63462 5480
rect 63314 5264 63370 5273
rect 63314 5199 63370 5208
rect 63512 4282 63540 6530
rect 63788 6526 63816 11886
rect 63776 6520 63828 6526
rect 63776 6462 63828 6468
rect 63880 6458 63908 12022
rect 63868 6452 63920 6458
rect 63868 6394 63920 6400
rect 63972 6361 64000 12158
rect 64064 6526 64092 45902
rect 64144 45756 64196 45762
rect 64144 45698 64196 45704
rect 64052 6520 64104 6526
rect 64052 6462 64104 6468
rect 63958 6352 64014 6361
rect 64156 6338 64184 45698
rect 64236 43852 64288 43858
rect 64236 43794 64288 43800
rect 64248 11218 64276 43794
rect 64420 31816 64472 31822
rect 64420 31758 64472 31764
rect 64328 29640 64380 29646
rect 64328 29582 64380 29588
rect 64236 11212 64288 11218
rect 64236 11154 64288 11160
rect 64236 11076 64288 11082
rect 64236 11018 64288 11024
rect 64248 7954 64276 11018
rect 64236 7948 64288 7954
rect 64236 7890 64288 7896
rect 64340 7546 64368 29582
rect 64328 7540 64380 7546
rect 64328 7482 64380 7488
rect 64328 6520 64380 6526
rect 64328 6462 64380 6468
rect 64236 6452 64288 6458
rect 64236 6394 64288 6400
rect 63958 6287 64014 6296
rect 64064 6310 64184 6338
rect 64064 6202 64092 6310
rect 63880 6174 64092 6202
rect 63880 5846 63908 6174
rect 64248 6066 64276 6394
rect 64340 6254 64368 6462
rect 64432 6390 64460 31758
rect 64512 27668 64564 27674
rect 64512 27610 64564 27616
rect 64420 6384 64472 6390
rect 64420 6326 64472 6332
rect 64328 6248 64380 6254
rect 64328 6190 64380 6196
rect 64524 6186 64552 27610
rect 64616 11354 64644 47330
rect 64972 44872 65024 44878
rect 64972 44814 65024 44820
rect 64880 41744 64932 41750
rect 64880 41686 64932 41692
rect 64892 39846 64920 41686
rect 64880 39840 64932 39846
rect 64880 39782 64932 39788
rect 64892 37398 64920 39782
rect 64880 37392 64932 37398
rect 64880 37334 64932 37340
rect 64892 35222 64920 37334
rect 64880 35216 64932 35222
rect 64880 35158 64932 35164
rect 64788 33992 64840 33998
rect 64788 33934 64840 33940
rect 64696 18760 64748 18766
rect 64696 18702 64748 18708
rect 64708 12481 64736 18702
rect 64694 12472 64750 12481
rect 64694 12407 64750 12416
rect 64696 12300 64748 12306
rect 64696 12242 64748 12248
rect 64604 11348 64656 11354
rect 64604 11290 64656 11296
rect 64604 11212 64656 11218
rect 64604 11154 64656 11160
rect 64512 6180 64564 6186
rect 64512 6122 64564 6128
rect 63972 6038 64276 6066
rect 63868 5840 63920 5846
rect 63868 5782 63920 5788
rect 63590 5264 63646 5273
rect 63590 5199 63646 5208
rect 63500 4276 63552 4282
rect 63500 4218 63552 4224
rect 63604 3097 63632 5199
rect 63972 3126 64000 6038
rect 64052 5772 64104 5778
rect 64052 5714 64104 5720
rect 64064 5642 64092 5714
rect 64052 5636 64104 5642
rect 64052 5578 64104 5584
rect 64188 5466 64540 5972
rect 64616 5778 64644 11154
rect 64708 7274 64736 12242
rect 64800 11506 64828 33934
rect 64892 33318 64920 35158
rect 64880 33312 64932 33318
rect 64880 33254 64932 33260
rect 64892 31142 64920 33254
rect 64880 31136 64932 31142
rect 64880 31078 64932 31084
rect 64892 28694 64920 31078
rect 64880 28688 64932 28694
rect 64880 28630 64932 28636
rect 64892 27062 64920 28630
rect 64880 27056 64932 27062
rect 64880 26998 64932 27004
rect 64984 23866 65012 44814
rect 64972 23860 65024 23866
rect 64972 23802 65024 23808
rect 64880 12776 64932 12782
rect 64880 12718 64932 12724
rect 64892 12434 64920 12718
rect 64892 12406 65012 12434
rect 64800 11478 64920 11506
rect 64788 11348 64840 11354
rect 64788 11290 64840 11296
rect 64696 7268 64748 7274
rect 64696 7210 64748 7216
rect 64604 5772 64656 5778
rect 64604 5714 64656 5720
rect 64800 5658 64828 11290
rect 64892 10606 64920 11478
rect 64880 10600 64932 10606
rect 64880 10542 64932 10548
rect 64880 10464 64932 10470
rect 64880 10406 64932 10412
rect 64892 6798 64920 10406
rect 64984 7818 65012 12406
rect 64972 7812 65024 7818
rect 64972 7754 65024 7760
rect 64970 7712 65026 7721
rect 64970 7647 65026 7656
rect 64880 6792 64932 6798
rect 64880 6734 64932 6740
rect 64984 6594 65012 7647
rect 64972 6588 65024 6594
rect 64972 6530 65024 6536
rect 64972 6248 65024 6254
rect 64972 6190 65024 6196
rect 64800 5630 64920 5658
rect 64788 5568 64840 5574
rect 64788 5510 64840 5516
rect 64188 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64540 5466
rect 64188 4588 64540 5414
rect 64188 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64540 4588
rect 64188 4508 64540 4532
rect 64188 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64540 4508
rect 64188 4428 64540 4452
rect 64188 4378 64216 4428
rect 64272 4378 64296 4428
rect 64352 4378 64376 4428
rect 64432 4378 64456 4428
rect 64512 4378 64540 4428
rect 64188 4326 64210 4378
rect 64272 4372 64274 4378
rect 64454 4372 64456 4378
rect 64262 4348 64274 4372
rect 64326 4348 64338 4372
rect 64390 4348 64402 4372
rect 64454 4348 64466 4372
rect 64272 4326 64274 4348
rect 64454 4326 64456 4348
rect 64518 4326 64540 4378
rect 64188 4292 64216 4326
rect 64272 4292 64296 4326
rect 64352 4292 64376 4326
rect 64432 4292 64456 4326
rect 64512 4292 64540 4326
rect 64188 3290 64540 4292
rect 64188 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64540 3290
rect 63960 3120 64012 3126
rect 63590 3088 63646 3097
rect 63224 3052 63276 3058
rect 63960 3062 64012 3068
rect 63590 3023 63646 3032
rect 63224 2994 63276 3000
rect 63040 2848 63092 2854
rect 63040 2790 63092 2796
rect 61836 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 62188 2746
rect 61836 2236 62188 2694
rect 62304 2440 62356 2446
rect 62304 2382 62356 2388
rect 61836 2180 61864 2236
rect 61920 2180 61944 2236
rect 62000 2180 62024 2236
rect 62080 2180 62104 2236
rect 62160 2180 62188 2236
rect 61836 2156 62188 2180
rect 61836 2100 61864 2156
rect 61920 2100 61944 2156
rect 62000 2100 62024 2156
rect 62080 2100 62104 2156
rect 62160 2100 62188 2156
rect 61836 2076 62188 2100
rect 61836 2020 61864 2076
rect 61920 2020 61944 2076
rect 62000 2020 62024 2076
rect 62080 2020 62104 2076
rect 62160 2020 62188 2076
rect 61836 1996 62188 2020
rect 61384 1964 61436 1970
rect 61384 1906 61436 1912
rect 61836 1940 61864 1996
rect 61920 1940 61944 1996
rect 62000 1940 62024 1996
rect 62080 1940 62104 1996
rect 62160 1940 62188 1996
rect 61108 1896 61160 1902
rect 61108 1838 61160 1844
rect 61016 1556 61068 1562
rect 61016 1498 61068 1504
rect 61120 800 61148 1838
rect 61836 1658 62188 1940
rect 61836 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 62188 1658
rect 61836 1040 62188 1606
rect 62316 1306 62344 2382
rect 62948 2304 63000 2310
rect 62948 2246 63000 2252
rect 62960 1970 62988 2246
rect 62948 1964 63000 1970
rect 62948 1906 63000 1912
rect 62396 1760 62448 1766
rect 62396 1702 62448 1708
rect 62408 1358 62436 1702
rect 62764 1420 62816 1426
rect 62764 1362 62816 1368
rect 62224 1278 62344 1306
rect 62396 1352 62448 1358
rect 62396 1294 62448 1300
rect 62224 800 62252 1278
rect 62776 800 62804 1362
rect 63052 1358 63080 2790
rect 63592 2372 63644 2378
rect 63592 2314 63644 2320
rect 63604 2106 63632 2314
rect 64188 2202 64540 3238
rect 64800 3058 64828 5510
rect 64892 5137 64920 5630
rect 64878 5128 64934 5137
rect 64878 5063 64934 5072
rect 64984 4078 65012 6190
rect 65076 5778 65104 71742
rect 65524 70032 65576 70038
rect 65524 69974 65576 69980
rect 65432 65680 65484 65686
rect 65432 65622 65484 65628
rect 65340 63572 65392 63578
rect 65340 63514 65392 63520
rect 65156 59152 65208 59158
rect 65156 59094 65208 59100
rect 65168 30938 65196 59094
rect 65248 49156 65300 49162
rect 65248 49098 65300 49104
rect 65260 44849 65288 49098
rect 65246 44840 65302 44849
rect 65246 44775 65302 44784
rect 65248 40996 65300 41002
rect 65248 40938 65300 40944
rect 65260 40905 65288 40938
rect 65246 40896 65302 40905
rect 65246 40831 65302 40840
rect 65248 38820 65300 38826
rect 65248 38762 65300 38768
rect 65260 38729 65288 38762
rect 65246 38720 65302 38729
rect 65246 38655 65302 38664
rect 65248 34536 65300 34542
rect 65248 34478 65300 34484
rect 65156 30932 65208 30938
rect 65156 30874 65208 30880
rect 65156 24336 65208 24342
rect 65156 24278 65208 24284
rect 65168 22166 65196 24278
rect 65156 22160 65208 22166
rect 65156 22102 65208 22108
rect 65168 20262 65196 22102
rect 65156 20256 65208 20262
rect 65156 20198 65208 20204
rect 65168 18018 65196 20198
rect 65156 18012 65208 18018
rect 65156 17954 65208 17960
rect 65168 15638 65196 17954
rect 65156 15632 65208 15638
rect 65156 15574 65208 15580
rect 65168 13734 65196 15574
rect 65156 13728 65208 13734
rect 65156 13670 65208 13676
rect 65168 11286 65196 13670
rect 65156 11280 65208 11286
rect 65156 11222 65208 11228
rect 65156 10600 65208 10606
rect 65156 10542 65208 10548
rect 65168 7070 65196 10542
rect 65156 7064 65208 7070
rect 65156 7006 65208 7012
rect 65156 6792 65208 6798
rect 65156 6734 65208 6740
rect 65064 5772 65116 5778
rect 65064 5714 65116 5720
rect 64972 4072 65024 4078
rect 64972 4014 65024 4020
rect 64788 3052 64840 3058
rect 64788 2994 64840 3000
rect 64604 2848 64656 2854
rect 64604 2790 64656 2796
rect 64188 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64540 2202
rect 63592 2100 63644 2106
rect 63592 2042 63644 2048
rect 63868 1896 63920 1902
rect 63868 1838 63920 1844
rect 63880 1562 63908 1838
rect 63868 1556 63920 1562
rect 63868 1498 63920 1504
rect 63040 1352 63092 1358
rect 63040 1294 63092 1300
rect 63868 1352 63920 1358
rect 63868 1294 63920 1300
rect 63880 800 63908 1294
rect 64188 1114 64540 2150
rect 64616 1970 64644 2790
rect 65168 2310 65196 6734
rect 65260 6497 65288 34478
rect 65352 33114 65380 63514
rect 65444 33658 65472 65622
rect 65536 36378 65564 69974
rect 65892 67856 65944 67862
rect 65892 67798 65944 67804
rect 65708 63232 65760 63238
rect 65708 63174 65760 63180
rect 65616 52488 65668 52494
rect 65616 52430 65668 52436
rect 65628 52154 65656 52430
rect 65616 52148 65668 52154
rect 65616 52090 65668 52096
rect 65524 36372 65576 36378
rect 65524 36314 65576 36320
rect 65616 33924 65668 33930
rect 65616 33866 65668 33872
rect 65432 33652 65484 33658
rect 65432 33594 65484 33600
rect 65628 33289 65656 33866
rect 65614 33280 65670 33289
rect 65614 33215 65670 33224
rect 65340 33108 65392 33114
rect 65340 33050 65392 33056
rect 65340 32224 65392 32230
rect 65340 32166 65392 32172
rect 65352 11370 65380 32166
rect 65432 30048 65484 30054
rect 65432 29990 65484 29996
rect 65444 11529 65472 29990
rect 65616 25696 65668 25702
rect 65616 25638 65668 25644
rect 65524 19168 65576 19174
rect 65522 19136 65524 19145
rect 65576 19136 65578 19145
rect 65522 19071 65578 19080
rect 65524 14816 65576 14822
rect 65524 14758 65576 14764
rect 65430 11520 65486 11529
rect 65430 11455 65486 11464
rect 65352 11342 65472 11370
rect 65340 11280 65392 11286
rect 65340 11222 65392 11228
rect 65352 9178 65380 11222
rect 65340 9172 65392 9178
rect 65340 9114 65392 9120
rect 65246 6488 65302 6497
rect 65246 6423 65302 6432
rect 65352 5302 65380 9114
rect 65444 5914 65472 11342
rect 65536 7342 65564 14758
rect 65524 7336 65576 7342
rect 65524 7278 65576 7284
rect 65524 6384 65576 6390
rect 65524 6326 65576 6332
rect 65432 5908 65484 5914
rect 65432 5850 65484 5856
rect 65340 5296 65392 5302
rect 65340 5238 65392 5244
rect 65536 2530 65564 6326
rect 65628 5166 65656 25638
rect 65720 7410 65748 63174
rect 65800 36576 65852 36582
rect 65800 36518 65852 36524
rect 65708 7404 65760 7410
rect 65708 7346 65760 7352
rect 65812 7018 65840 36518
rect 65904 35290 65932 67798
rect 66076 61328 66128 61334
rect 66076 61270 66128 61276
rect 65984 54528 66036 54534
rect 65984 54470 66036 54476
rect 65892 35284 65944 35290
rect 65892 35226 65944 35232
rect 65892 27872 65944 27878
rect 65892 27814 65944 27820
rect 65720 6990 65840 7018
rect 65720 6633 65748 6990
rect 65800 6860 65852 6866
rect 65800 6802 65852 6808
rect 65706 6624 65762 6633
rect 65706 6559 65762 6568
rect 65616 5160 65668 5166
rect 65616 5102 65668 5108
rect 65444 2502 65564 2530
rect 65812 2514 65840 6802
rect 65904 5370 65932 27814
rect 65996 5817 66024 54470
rect 66088 32026 66116 61270
rect 66076 32020 66128 32026
rect 66076 31962 66128 31968
rect 66076 23520 66128 23526
rect 66076 23462 66128 23468
rect 65982 5808 66038 5817
rect 65982 5743 66038 5752
rect 65892 5364 65944 5370
rect 65892 5306 65944 5312
rect 66088 5098 66116 23462
rect 66180 5778 66208 74054
rect 66272 39642 66300 76502
rect 66352 51536 66404 51542
rect 66352 51478 66404 51484
rect 66260 39636 66312 39642
rect 66260 39578 66312 39584
rect 66260 28552 66312 28558
rect 66260 28494 66312 28500
rect 66168 5772 66220 5778
rect 66168 5714 66220 5720
rect 66076 5092 66128 5098
rect 66076 5034 66128 5040
rect 66272 3670 66300 28494
rect 66364 26926 66392 51478
rect 66456 40730 66484 78678
rect 66628 72208 66680 72214
rect 66628 72150 66680 72156
rect 66536 68944 66588 68950
rect 66536 68886 66588 68892
rect 66444 40724 66496 40730
rect 66444 40666 66496 40672
rect 66548 35766 66576 68886
rect 66640 37194 66668 72150
rect 66904 53168 66956 53174
rect 66904 53110 66956 53116
rect 66812 52624 66864 52630
rect 66812 52566 66864 52572
rect 66628 37188 66680 37194
rect 66628 37130 66680 37136
rect 66824 35894 66852 52566
rect 66732 35866 66852 35894
rect 66536 35760 66588 35766
rect 66536 35702 66588 35708
rect 66732 35170 66760 35866
rect 66548 35142 66760 35170
rect 66444 33040 66496 33046
rect 66444 32982 66496 32988
rect 66456 29850 66484 32982
rect 66444 29844 66496 29850
rect 66444 29786 66496 29792
rect 66444 29640 66496 29646
rect 66444 29582 66496 29588
rect 66352 26920 66404 26926
rect 66352 26862 66404 26868
rect 66352 24200 66404 24206
rect 66352 24142 66404 24148
rect 66364 23497 66392 24142
rect 66350 23488 66406 23497
rect 66350 23423 66406 23432
rect 66350 23352 66406 23361
rect 66350 23287 66406 23296
rect 66260 3664 66312 3670
rect 66260 3606 66312 3612
rect 66364 3602 66392 23287
rect 66456 6458 66484 29582
rect 66548 27606 66576 35142
rect 66628 35080 66680 35086
rect 66628 35022 66680 35028
rect 66536 27600 66588 27606
rect 66536 27542 66588 27548
rect 66536 26376 66588 26382
rect 66536 26318 66588 26324
rect 66548 23798 66576 26318
rect 66536 23792 66588 23798
rect 66536 23734 66588 23740
rect 66536 23656 66588 23662
rect 66536 23598 66588 23604
rect 66548 23497 66576 23598
rect 66534 23488 66590 23497
rect 66534 23423 66590 23432
rect 66536 23112 66588 23118
rect 66536 23054 66588 23060
rect 66444 6452 66496 6458
rect 66444 6394 66496 6400
rect 66548 6254 66576 23054
rect 66640 6866 66668 35022
rect 66916 34202 66944 53110
rect 67008 42770 67036 83098
rect 69664 83020 69716 83026
rect 69664 82962 69716 82968
rect 67088 80980 67140 80986
rect 67088 80922 67140 80928
rect 66996 42764 67048 42770
rect 66996 42706 67048 42712
rect 67100 41818 67128 80922
rect 68468 76492 68520 76498
rect 68468 76434 68520 76440
rect 67824 74656 67876 74662
rect 67824 74598 67876 74604
rect 67548 56976 67600 56982
rect 67548 56918 67600 56924
rect 67180 46980 67232 46986
rect 67180 46922 67232 46928
rect 67088 41812 67140 41818
rect 67088 41754 67140 41760
rect 66996 38344 67048 38350
rect 66996 38286 67048 38292
rect 66904 34196 66956 34202
rect 66904 34138 66956 34144
rect 66720 33448 66772 33454
rect 66720 33390 66772 33396
rect 66628 6860 66680 6866
rect 66628 6802 66680 6808
rect 66732 6390 66760 33390
rect 67008 31090 67036 38286
rect 67088 31816 67140 31822
rect 67088 31758 67140 31764
rect 66916 31062 67036 31090
rect 66812 30728 66864 30734
rect 66812 30670 66864 30676
rect 66824 6798 66852 30670
rect 66812 6792 66864 6798
rect 66812 6734 66864 6740
rect 66720 6384 66772 6390
rect 66720 6326 66772 6332
rect 66536 6248 66588 6254
rect 66536 6190 66588 6196
rect 66444 5568 66496 5574
rect 66444 5510 66496 5516
rect 66352 3596 66404 3602
rect 66352 3538 66404 3544
rect 66456 3058 66484 5510
rect 66444 3052 66496 3058
rect 66444 2994 66496 3000
rect 66260 2848 66312 2854
rect 66260 2790 66312 2796
rect 65800 2508 65852 2514
rect 65156 2304 65208 2310
rect 65156 2246 65208 2252
rect 64604 1964 64656 1970
rect 64604 1906 64656 1912
rect 64696 1896 64748 1902
rect 64696 1838 64748 1844
rect 64188 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64540 1114
rect 64188 1040 64540 1062
rect 64432 870 64552 898
rect 64432 800 64460 870
rect 44652 734 44864 762
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64524 762 64552 870
rect 64708 762 64736 1838
rect 65444 1834 65472 2502
rect 65800 2450 65852 2456
rect 65524 2440 65576 2446
rect 65524 2382 65576 2388
rect 65432 1828 65484 1834
rect 65432 1770 65484 1776
rect 65156 1760 65208 1766
rect 65156 1702 65208 1708
rect 65168 1358 65196 1702
rect 65156 1352 65208 1358
rect 65156 1294 65208 1300
rect 65536 800 65564 2382
rect 66076 2304 66128 2310
rect 66076 2246 66128 2252
rect 66088 1970 66116 2246
rect 66076 1964 66128 1970
rect 66076 1906 66128 1912
rect 66272 1358 66300 2790
rect 66916 2038 66944 31062
rect 66996 27464 67048 27470
rect 66996 27406 67048 27412
rect 67008 23905 67036 27406
rect 66994 23896 67050 23905
rect 66994 23831 67050 23840
rect 66996 23792 67048 23798
rect 66996 23734 67048 23740
rect 67008 3466 67036 23734
rect 67100 3534 67128 31758
rect 67192 11082 67220 46922
rect 67456 39432 67508 39438
rect 67456 39374 67508 39380
rect 67272 37256 67324 37262
rect 67272 37198 67324 37204
rect 67180 11076 67232 11082
rect 67180 11018 67232 11024
rect 67088 3528 67140 3534
rect 67088 3470 67140 3476
rect 66996 3460 67048 3466
rect 66996 3402 67048 3408
rect 67284 2530 67312 37198
rect 67364 36168 67416 36174
rect 67364 36110 67416 36116
rect 67376 2650 67404 36110
rect 67364 2644 67416 2650
rect 67364 2586 67416 2592
rect 67284 2502 67404 2530
rect 67468 2514 67496 39374
rect 67560 33046 67588 56918
rect 67732 54868 67784 54874
rect 67732 54810 67784 54816
rect 67640 50516 67692 50522
rect 67640 50458 67692 50464
rect 67548 33040 67600 33046
rect 67548 32982 67600 32988
rect 67548 32904 67600 32910
rect 67548 32846 67600 32852
rect 67560 4146 67588 32846
rect 67652 26586 67680 50458
rect 67744 28762 67772 54810
rect 67836 38554 67864 74598
rect 68376 47048 68428 47054
rect 68376 46990 68428 46996
rect 68192 44532 68244 44538
rect 68192 44474 68244 44480
rect 67916 38752 67968 38758
rect 67916 38694 67968 38700
rect 67824 38548 67876 38554
rect 67824 38490 67876 38496
rect 67732 28756 67784 28762
rect 67732 28698 67784 28704
rect 67640 26580 67692 26586
rect 67640 26522 67692 26528
rect 67824 21140 67876 21146
rect 67824 21082 67876 21088
rect 67640 14612 67692 14618
rect 67640 14554 67692 14560
rect 67652 5846 67680 14554
rect 67732 12640 67784 12646
rect 67732 12582 67784 12588
rect 67744 6118 67772 12582
rect 67836 6322 67864 21082
rect 67824 6316 67876 6322
rect 67824 6258 67876 6264
rect 67732 6112 67784 6118
rect 67732 6054 67784 6060
rect 67640 5840 67692 5846
rect 67640 5782 67692 5788
rect 67928 4622 67956 38694
rect 68100 36304 68152 36310
rect 68100 36246 68152 36252
rect 68008 35692 68060 35698
rect 68008 35634 68060 35640
rect 67916 4616 67968 4622
rect 67916 4558 67968 4564
rect 67548 4140 67600 4146
rect 67548 4082 67600 4088
rect 68020 2774 68048 35634
rect 68112 16574 68140 36246
rect 68204 23322 68232 44474
rect 68284 44464 68336 44470
rect 68284 44406 68336 44412
rect 68296 24410 68324 44406
rect 68284 24404 68336 24410
rect 68284 24346 68336 24352
rect 68192 23316 68244 23322
rect 68192 23258 68244 23264
rect 68112 16546 68232 16574
rect 68100 5568 68152 5574
rect 68100 5510 68152 5516
rect 68112 3058 68140 5510
rect 68204 5030 68232 16546
rect 68388 7478 68416 46990
rect 68376 7472 68428 7478
rect 68376 7414 68428 7420
rect 68480 5778 68508 76434
rect 69020 59084 69072 59090
rect 69020 59026 69072 59032
rect 68560 43104 68612 43110
rect 68560 43046 68612 43052
rect 68468 5772 68520 5778
rect 68468 5714 68520 5720
rect 68192 5024 68244 5030
rect 68192 4966 68244 4972
rect 68572 4486 68600 43046
rect 68652 40928 68704 40934
rect 68652 40870 68704 40876
rect 68664 4554 68692 40870
rect 68836 27056 68888 27062
rect 68836 26998 68888 27004
rect 68744 26988 68796 26994
rect 68744 26930 68796 26936
rect 68652 4548 68704 4554
rect 68652 4490 68704 4496
rect 68560 4480 68612 4486
rect 68560 4422 68612 4428
rect 68100 3052 68152 3058
rect 68100 2994 68152 3000
rect 68284 2848 68336 2854
rect 68284 2790 68336 2796
rect 67928 2746 68048 2774
rect 67272 2440 67324 2446
rect 67272 2382 67324 2388
rect 67284 2106 67312 2382
rect 67272 2100 67324 2106
rect 67272 2042 67324 2048
rect 66904 2032 66956 2038
rect 66904 1974 66956 1980
rect 67180 1964 67232 1970
rect 67180 1906 67232 1912
rect 66260 1352 66312 1358
rect 66260 1294 66312 1300
rect 66076 1284 66128 1290
rect 66076 1226 66128 1232
rect 66088 800 66116 1226
rect 67192 800 67220 1906
rect 67376 1222 67404 2502
rect 67456 2508 67508 2514
rect 67456 2450 67508 2456
rect 67928 2038 67956 2746
rect 67916 2032 67968 2038
rect 67916 1974 67968 1980
rect 67732 1420 67784 1426
rect 67732 1362 67784 1368
rect 67364 1216 67416 1222
rect 67364 1158 67416 1164
rect 67744 800 67772 1362
rect 68296 1358 68324 2790
rect 68756 2582 68784 26930
rect 68848 5642 68876 26998
rect 68928 23248 68980 23254
rect 68928 23190 68980 23196
rect 68940 6866 68968 23190
rect 68928 6860 68980 6866
rect 68928 6802 68980 6808
rect 68836 5636 68888 5642
rect 68836 5578 68888 5584
rect 69032 4690 69060 59026
rect 69204 40520 69256 40526
rect 69204 40462 69256 40468
rect 69020 4684 69072 4690
rect 69020 4626 69072 4632
rect 68744 2576 68796 2582
rect 68744 2518 68796 2524
rect 69216 2038 69244 40462
rect 69676 5302 69704 82962
rect 71836 82236 72188 83206
rect 71836 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 72188 82236
rect 71836 82170 72188 82180
rect 71836 82118 71858 82170
rect 71910 82156 71922 82170
rect 71974 82156 71986 82170
rect 72038 82156 72050 82170
rect 72102 82156 72114 82170
rect 71920 82118 71922 82156
rect 72102 82118 72104 82156
rect 72166 82118 72188 82170
rect 71836 82100 71864 82118
rect 71920 82100 71944 82118
rect 72000 82100 72024 82118
rect 72080 82100 72104 82118
rect 72160 82100 72188 82118
rect 71836 82076 72188 82100
rect 71836 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 72188 82076
rect 71836 81996 72188 82020
rect 71836 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 72188 81996
rect 71836 81082 72188 81940
rect 71836 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 72188 81082
rect 69756 80844 69808 80850
rect 69756 80786 69808 80792
rect 69664 5296 69716 5302
rect 69664 5238 69716 5244
rect 69768 5098 69796 80786
rect 71836 79994 72188 81030
rect 71836 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 72188 79994
rect 71836 78906 72188 79942
rect 71836 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 72188 78906
rect 69940 78668 69992 78674
rect 69940 78610 69992 78616
rect 69952 5166 69980 78610
rect 71836 77818 72188 78854
rect 71836 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 72188 77818
rect 71836 76730 72188 77766
rect 71836 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 72188 76730
rect 71836 75642 72188 76678
rect 71836 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 72188 75642
rect 71836 74554 72188 75590
rect 71836 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 72188 74554
rect 71836 73466 72188 74502
rect 71836 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 72188 73466
rect 71836 72378 72188 73414
rect 71836 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 72188 72378
rect 71836 72236 72188 72326
rect 71836 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 72188 72236
rect 71836 72156 72188 72180
rect 71836 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 72188 72156
rect 71836 72076 72188 72100
rect 71836 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 72188 72076
rect 71836 71996 72188 72020
rect 71836 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 72188 71996
rect 71836 71290 72188 71940
rect 71836 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 72188 71290
rect 71836 70202 72188 71238
rect 71836 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 72188 70202
rect 71836 69114 72188 70150
rect 71836 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 72188 69114
rect 71836 68026 72188 69062
rect 71836 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 72188 68026
rect 71836 66938 72188 67974
rect 71836 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 72188 66938
rect 71836 65850 72188 66886
rect 71836 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 72188 65850
rect 70400 65612 70452 65618
rect 70400 65554 70452 65560
rect 70032 42696 70084 42702
rect 70032 42638 70084 42644
rect 69940 5160 69992 5166
rect 69940 5102 69992 5108
rect 69756 5092 69808 5098
rect 69756 5034 69808 5040
rect 69848 5024 69900 5030
rect 69848 4966 69900 4972
rect 69860 3058 69888 4966
rect 69848 3052 69900 3058
rect 69848 2994 69900 3000
rect 69664 2848 69716 2854
rect 69664 2790 69716 2796
rect 69388 2304 69440 2310
rect 69388 2246 69440 2252
rect 69204 2032 69256 2038
rect 69204 1974 69256 1980
rect 69400 1970 69428 2246
rect 69676 1970 69704 2790
rect 69940 2440 69992 2446
rect 69940 2382 69992 2388
rect 69388 1964 69440 1970
rect 69388 1906 69440 1912
rect 69664 1964 69716 1970
rect 69664 1906 69716 1912
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 68284 1352 68336 1358
rect 68284 1294 68336 1300
rect 68836 1352 68888 1358
rect 68836 1294 68888 1300
rect 68848 800 68876 1294
rect 69400 800 69428 1770
rect 69952 1562 69980 2382
rect 69940 1556 69992 1562
rect 69940 1498 69992 1504
rect 70044 1290 70072 42638
rect 70124 41608 70176 41614
rect 70124 41550 70176 41556
rect 70136 2038 70164 41550
rect 70412 6089 70440 65554
rect 71836 64762 72188 65798
rect 71836 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 72188 64762
rect 71836 63674 72188 64710
rect 71836 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 72188 63674
rect 71836 62586 72188 63622
rect 71836 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 72188 62586
rect 71836 62236 72188 62534
rect 71836 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 72188 62236
rect 71836 62156 72188 62180
rect 71836 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 72188 62156
rect 71836 62076 72188 62100
rect 71836 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 72188 62076
rect 71836 61996 72188 62020
rect 71836 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 72188 61996
rect 71836 61498 72188 61940
rect 71836 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 72188 61498
rect 71836 60410 72188 61446
rect 71836 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 72188 60410
rect 71836 59322 72188 60358
rect 71836 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 72188 59322
rect 71836 58234 72188 59270
rect 71836 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 72188 58234
rect 71836 57146 72188 58182
rect 71836 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 72188 57146
rect 70492 56908 70544 56914
rect 70492 56850 70544 56856
rect 70398 6080 70454 6089
rect 70398 6015 70454 6024
rect 70504 4214 70532 56850
rect 71836 56058 72188 57094
rect 71836 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 72188 56058
rect 71836 54970 72188 56006
rect 71836 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 72188 54970
rect 71836 53882 72188 54918
rect 71836 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 72188 53882
rect 71836 52794 72188 53830
rect 71836 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 72188 52794
rect 71836 52236 72188 52742
rect 71836 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 72188 52236
rect 71836 52156 72188 52180
rect 71836 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 72188 52156
rect 71836 52076 72188 52100
rect 71836 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 72188 52076
rect 71836 51996 72188 52020
rect 71836 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 72188 51996
rect 71836 51706 72188 51940
rect 71836 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 72188 51706
rect 71836 50618 72188 51654
rect 71836 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 72188 50618
rect 71836 49530 72188 50566
rect 71836 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 72188 49530
rect 71836 48442 72188 49478
rect 71836 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 72188 48442
rect 71836 47354 72188 48390
rect 71836 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 72188 47354
rect 71836 46266 72188 47302
rect 71836 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 72188 46266
rect 71836 45178 72188 46214
rect 71836 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 72188 45178
rect 71836 44090 72188 45126
rect 71836 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 72188 44090
rect 71836 43002 72188 44038
rect 71836 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 72188 43002
rect 71836 42236 72188 42950
rect 71836 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 72188 42236
rect 71836 42156 72188 42180
rect 71836 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 72188 42156
rect 71836 42076 72188 42100
rect 71836 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 72188 42076
rect 71836 41996 72188 42020
rect 71836 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 72188 41996
rect 71836 41914 72188 41940
rect 71836 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 72188 41914
rect 71836 40826 72188 41862
rect 71836 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 72188 40826
rect 71836 39738 72188 40774
rect 71836 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 72188 39738
rect 71836 38650 72188 39686
rect 71836 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 72188 38650
rect 71836 37562 72188 38598
rect 71836 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 72188 37562
rect 71836 36474 72188 37510
rect 71836 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 72188 36474
rect 71836 35386 72188 36422
rect 71836 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 72188 35386
rect 71836 34298 72188 35334
rect 71836 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 72188 34298
rect 71836 33210 72188 34246
rect 71836 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 72188 33210
rect 71836 32236 72188 33158
rect 71836 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 72188 32236
rect 71836 32156 72188 32180
rect 71836 32122 71864 32156
rect 71920 32122 71944 32156
rect 72000 32122 72024 32156
rect 72080 32122 72104 32156
rect 72160 32122 72188 32156
rect 71836 32070 71858 32122
rect 71920 32100 71922 32122
rect 72102 32100 72104 32122
rect 71910 32076 71922 32100
rect 71974 32076 71986 32100
rect 72038 32076 72050 32100
rect 72102 32076 72114 32100
rect 71920 32070 71922 32076
rect 72102 32070 72104 32076
rect 72166 32070 72188 32122
rect 71836 32020 71864 32070
rect 71920 32020 71944 32070
rect 72000 32020 72024 32070
rect 72080 32020 72104 32070
rect 72160 32020 72188 32070
rect 71836 31996 72188 32020
rect 71836 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 72188 31996
rect 71836 31034 72188 31940
rect 71836 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 72188 31034
rect 71836 29946 72188 30982
rect 71836 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 72188 29946
rect 71836 28858 72188 29894
rect 71836 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 72188 28858
rect 71836 27770 72188 28806
rect 71836 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 72188 27770
rect 71836 26682 72188 27718
rect 71836 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 72188 26682
rect 71836 25594 72188 26630
rect 71836 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 72188 25594
rect 71836 24506 72188 25542
rect 71836 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 72188 24506
rect 71836 23418 72188 24454
rect 71836 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 72188 23418
rect 71836 22330 72188 23366
rect 71836 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 72188 22330
rect 71836 22236 72188 22278
rect 71836 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 72188 22236
rect 71836 22156 72188 22180
rect 71836 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 72188 22156
rect 71836 22076 72188 22100
rect 71836 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 72188 22076
rect 71836 21996 72188 22020
rect 71836 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 72188 21996
rect 70584 21548 70636 21554
rect 70584 21490 70636 21496
rect 70596 6662 70624 21490
rect 71836 21242 72188 21940
rect 71836 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 72188 21242
rect 71836 20154 72188 21190
rect 71836 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 72188 20154
rect 71836 19066 72188 20102
rect 71836 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 72188 19066
rect 71836 17978 72188 19014
rect 71836 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 72188 17978
rect 70676 17196 70728 17202
rect 70676 17138 70728 17144
rect 70688 6730 70716 17138
rect 71836 16890 72188 17926
rect 71836 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 72188 16890
rect 71836 15802 72188 16838
rect 71836 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 72188 15802
rect 71836 14714 72188 15750
rect 71836 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 72188 14714
rect 71836 13626 72188 14662
rect 71836 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 72188 13626
rect 71836 12538 72188 13574
rect 71836 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 72188 12538
rect 71836 12236 72188 12486
rect 71836 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 72188 12236
rect 71836 12156 72188 12180
rect 71836 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 72188 12156
rect 71836 12076 72188 12100
rect 71836 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 72188 12076
rect 71836 11996 72188 12020
rect 71836 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 72188 11996
rect 71836 11450 72188 11940
rect 71836 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 72188 11450
rect 71836 10362 72188 11398
rect 71836 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 72188 10362
rect 71836 9274 72188 10310
rect 71836 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 72188 9274
rect 71836 8186 72188 9222
rect 71836 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 72188 8186
rect 71836 7098 72188 8134
rect 71836 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 72188 7098
rect 70676 6724 70728 6730
rect 70676 6666 70728 6672
rect 70584 6656 70636 6662
rect 70584 6598 70636 6604
rect 71836 6010 72188 7046
rect 71836 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 72188 6010
rect 71412 5024 71464 5030
rect 71412 4966 71464 4972
rect 70492 4208 70544 4214
rect 70492 4150 70544 4156
rect 71424 3058 71452 4966
rect 71836 4922 72188 5958
rect 74188 85978 74540 86000
rect 74188 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74540 85978
rect 74188 84890 74540 85926
rect 74188 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74540 84890
rect 74188 84588 74540 84838
rect 74188 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 74540 84588
rect 74188 84508 74540 84532
rect 74188 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 74540 84508
rect 74188 84428 74540 84452
rect 74188 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 74540 84428
rect 74188 84348 74540 84372
rect 74188 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 74540 84348
rect 74188 83802 74540 84292
rect 74188 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74540 83802
rect 74188 82714 74540 83750
rect 74188 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74540 82714
rect 74188 81626 74540 82662
rect 74188 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74540 81626
rect 74188 80538 74540 81574
rect 74188 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74540 80538
rect 74188 79450 74540 80486
rect 74188 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74540 79450
rect 74188 78362 74540 79398
rect 74188 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74540 78362
rect 74188 77274 74540 78310
rect 74188 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74540 77274
rect 74188 76186 74540 77222
rect 74188 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74540 76186
rect 74188 75098 74540 76134
rect 74188 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74540 75098
rect 74188 74588 74540 75046
rect 74188 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 74540 74588
rect 74188 74508 74540 74532
rect 74188 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 74540 74508
rect 74188 74428 74540 74452
rect 74188 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 74540 74428
rect 74188 74348 74540 74372
rect 74188 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 74540 74348
rect 74188 74010 74540 74292
rect 74188 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74540 74010
rect 74188 72922 74540 73958
rect 74188 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74540 72922
rect 74188 71834 74540 72870
rect 74188 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74540 71834
rect 74188 70746 74540 71782
rect 74188 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74540 70746
rect 74188 69658 74540 70694
rect 74188 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74540 69658
rect 74188 68570 74540 69606
rect 74188 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74540 68570
rect 74188 67482 74540 68518
rect 74188 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74540 67482
rect 74188 66394 74540 67430
rect 74188 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74540 66394
rect 74188 65306 74540 66342
rect 74188 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74540 65306
rect 74188 64588 74540 65254
rect 74188 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 74540 64588
rect 74188 64508 74540 64532
rect 74188 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 74540 64508
rect 74188 64428 74540 64452
rect 74188 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 74540 64428
rect 74188 64348 74540 64372
rect 74188 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 74540 64348
rect 74188 64218 74540 64292
rect 74188 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74540 64218
rect 74188 63130 74540 64166
rect 74188 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74540 63130
rect 74188 62042 74540 63078
rect 74188 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74540 62042
rect 74188 60954 74540 61990
rect 74188 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74540 60954
rect 74188 59866 74540 60902
rect 74188 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74540 59866
rect 74188 58778 74540 59814
rect 74188 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74540 58778
rect 74188 57690 74540 58726
rect 74188 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74540 57690
rect 74188 56602 74540 57638
rect 74188 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74540 56602
rect 74188 55514 74540 56550
rect 74188 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74540 55514
rect 74188 54588 74540 55462
rect 74188 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 74540 54588
rect 74188 54508 74540 54532
rect 74188 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 74540 54508
rect 74188 54428 74540 54452
rect 74188 54426 74216 54428
rect 74272 54426 74296 54428
rect 74352 54426 74376 54428
rect 74432 54426 74456 54428
rect 74512 54426 74540 54428
rect 74188 54374 74210 54426
rect 74272 54374 74274 54426
rect 74454 54374 74456 54426
rect 74518 54374 74540 54426
rect 74188 54372 74216 54374
rect 74272 54372 74296 54374
rect 74352 54372 74376 54374
rect 74432 54372 74456 54374
rect 74512 54372 74540 54374
rect 74188 54348 74540 54372
rect 74188 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 74540 54348
rect 74188 53338 74540 54292
rect 74188 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74540 53338
rect 74188 52250 74540 53286
rect 74188 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74540 52250
rect 74188 51162 74540 52198
rect 74188 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74540 51162
rect 74188 50074 74540 51110
rect 74188 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74540 50074
rect 74188 48986 74540 50022
rect 74188 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74540 48986
rect 74188 47898 74540 48934
rect 74188 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74540 47898
rect 74188 46810 74540 47846
rect 74188 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74540 46810
rect 74188 45722 74540 46758
rect 74188 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74540 45722
rect 74188 44634 74540 45670
rect 74188 44582 74210 44634
rect 74262 44588 74274 44634
rect 74326 44588 74338 44634
rect 74390 44588 74402 44634
rect 74454 44588 74466 44634
rect 74272 44582 74274 44588
rect 74454 44582 74456 44588
rect 74518 44582 74540 44634
rect 74188 44532 74216 44582
rect 74272 44532 74296 44582
rect 74352 44532 74376 44582
rect 74432 44532 74456 44582
rect 74512 44532 74540 44582
rect 74188 44508 74540 44532
rect 74188 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 74540 44508
rect 74188 44428 74540 44452
rect 74188 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 74540 44428
rect 74188 44348 74540 44372
rect 74188 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 74540 44348
rect 74188 43546 74540 44292
rect 74188 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74540 43546
rect 74188 42458 74540 43494
rect 74188 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74540 42458
rect 74188 41370 74540 42406
rect 74188 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74540 41370
rect 74188 40282 74540 41318
rect 74188 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74540 40282
rect 74188 39194 74540 40230
rect 74188 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74540 39194
rect 74188 38106 74540 39142
rect 74188 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74540 38106
rect 74188 37018 74540 38054
rect 74188 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74540 37018
rect 74188 35930 74540 36966
rect 74188 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74540 35930
rect 74188 34842 74540 35878
rect 74188 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74540 34842
rect 74188 34588 74540 34790
rect 74188 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 74540 34588
rect 74188 34508 74540 34532
rect 74188 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 74540 34508
rect 74188 34428 74540 34452
rect 74188 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 74540 34428
rect 74188 34348 74540 34372
rect 74188 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 74540 34348
rect 74188 33754 74540 34292
rect 74188 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74540 33754
rect 74188 32666 74540 33702
rect 74188 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74540 32666
rect 74188 31578 74540 32614
rect 74188 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74540 31578
rect 74188 30490 74540 31526
rect 74188 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74540 30490
rect 74188 29402 74540 30438
rect 74188 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74540 29402
rect 74188 28314 74540 29350
rect 74188 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74540 28314
rect 74188 27226 74540 28262
rect 74188 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74540 27226
rect 74188 26138 74540 27174
rect 74188 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74540 26138
rect 74188 25050 74540 26086
rect 74188 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74540 25050
rect 74188 24588 74540 24998
rect 74188 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 74540 24588
rect 74188 24508 74540 24532
rect 74188 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 74540 24508
rect 74188 24428 74540 24452
rect 74188 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 74540 24428
rect 74188 24348 74540 24372
rect 74188 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 74540 24348
rect 74188 23962 74540 24292
rect 74188 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74540 23962
rect 74188 22874 74540 23910
rect 74188 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74540 22874
rect 74188 21786 74540 22822
rect 74188 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74540 21786
rect 74188 20698 74540 21734
rect 74188 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74540 20698
rect 74188 19610 74540 20646
rect 74188 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74540 19610
rect 74188 18522 74540 19558
rect 74188 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74540 18522
rect 74188 17434 74540 18470
rect 74188 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74540 17434
rect 74188 16346 74540 17382
rect 74188 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74540 16346
rect 74188 15258 74540 16294
rect 74188 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74540 15258
rect 74188 14588 74540 15206
rect 74188 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 74540 14588
rect 74188 14508 74540 14532
rect 74188 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 74540 14508
rect 74188 14428 74540 14452
rect 74188 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 74540 14428
rect 74188 14348 74540 14372
rect 74188 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 74540 14348
rect 74188 14170 74540 14292
rect 74188 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74540 14170
rect 74188 13082 74540 14118
rect 74188 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74540 13082
rect 74188 11994 74540 13030
rect 74188 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74540 11994
rect 74188 10906 74540 11942
rect 74188 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74540 10906
rect 74188 9818 74540 10854
rect 74188 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74540 9818
rect 74188 8730 74540 9766
rect 74188 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74540 8730
rect 74188 7642 74540 8678
rect 74188 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74540 7642
rect 74188 6554 74540 7590
rect 74188 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74540 6554
rect 74188 5466 74540 6502
rect 74188 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74540 5466
rect 73252 5024 73304 5030
rect 73252 4966 73304 4972
rect 71836 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 72188 4922
rect 71836 3834 72188 4870
rect 71836 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 72188 3834
rect 71412 3052 71464 3058
rect 71412 2994 71464 3000
rect 71228 2848 71280 2854
rect 71228 2790 71280 2796
rect 70492 2440 70544 2446
rect 70492 2382 70544 2388
rect 70124 2032 70176 2038
rect 70124 1974 70176 1980
rect 70032 1284 70084 1290
rect 70032 1226 70084 1232
rect 70504 800 70532 2382
rect 71044 2304 71096 2310
rect 71044 2246 71096 2252
rect 71056 1970 71084 2246
rect 71044 1964 71096 1970
rect 71044 1906 71096 1912
rect 71044 1420 71096 1426
rect 71044 1362 71096 1368
rect 71056 800 71084 1362
rect 71240 1358 71268 2790
rect 71836 2746 72188 3782
rect 73264 3058 73292 4966
rect 74188 4588 74540 5414
rect 74188 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 74540 4588
rect 74188 4508 74540 4532
rect 74188 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 74540 4508
rect 74188 4428 74540 4452
rect 74188 4378 74216 4428
rect 74272 4378 74296 4428
rect 74352 4378 74376 4428
rect 74432 4378 74456 4428
rect 74512 4378 74540 4428
rect 74188 4326 74210 4378
rect 74272 4372 74274 4378
rect 74454 4372 74456 4378
rect 74262 4348 74274 4372
rect 74326 4348 74338 4372
rect 74390 4348 74402 4372
rect 74454 4348 74466 4372
rect 74272 4326 74274 4348
rect 74454 4326 74456 4348
rect 74518 4326 74540 4378
rect 74188 4292 74216 4326
rect 74272 4292 74296 4326
rect 74352 4292 74376 4326
rect 74432 4292 74456 4326
rect 74512 4292 74540 4326
rect 74188 3290 74540 4292
rect 74188 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74540 3290
rect 73252 3052 73304 3058
rect 73252 2994 73304 3000
rect 73252 2848 73304 2854
rect 73252 2790 73304 2796
rect 71836 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 72188 2746
rect 71836 2236 72188 2694
rect 71836 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 72188 2236
rect 71836 2156 72188 2180
rect 71836 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 72188 2156
rect 71836 2076 72188 2100
rect 71836 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 72188 2076
rect 71836 1996 72188 2020
rect 71836 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 72188 1996
rect 71836 1658 72188 1940
rect 72240 1896 72292 1902
rect 72240 1838 72292 1844
rect 71836 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 72188 1658
rect 71228 1352 71280 1358
rect 71228 1294 71280 1300
rect 71836 1040 72188 1606
rect 72252 898 72280 1838
rect 73160 1760 73212 1766
rect 73160 1702 73212 1708
rect 73172 1358 73200 1702
rect 73264 1358 73292 2790
rect 74188 2202 74540 3238
rect 74188 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74540 2202
rect 73160 1352 73212 1358
rect 73160 1294 73212 1300
rect 73252 1352 73304 1358
rect 73252 1294 73304 1300
rect 72700 1216 72752 1222
rect 72700 1158 72752 1164
rect 72160 870 72280 898
rect 72160 800 72188 870
rect 72712 800 72740 1158
rect 74188 1114 74540 2150
rect 74188 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74540 1114
rect 74188 1040 74540 1062
rect 64524 734 64736 762
rect 64970 0 65026 800
rect 65522 0 65578 800
rect 66074 0 66130 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68282 0 68338 800
rect 68834 0 68890 800
rect 69386 0 69442 800
rect 69938 0 69994 800
rect 70490 0 70546 800
rect 71042 0 71098 800
rect 71594 0 71650 800
rect 72146 0 72202 800
rect 72698 0 72754 800
<< via2 >>
rect 2044 84532 2100 84588
rect 2044 84452 2100 84508
rect 2044 84372 2100 84428
rect 2044 84292 2100 84348
rect 5540 84532 5596 84588
rect 5540 84452 5596 84508
rect 5540 84372 5596 84428
rect 5540 84292 5596 84348
rect 8430 84532 8486 84588
rect 8430 84452 8486 84508
rect 8430 84372 8486 84428
rect 8430 84292 8486 84348
rect 11320 84532 11376 84588
rect 11320 84452 11376 84508
rect 11320 84372 11376 84428
rect 11320 84292 11376 84348
rect 14210 84532 14266 84588
rect 14210 84452 14266 84508
rect 14210 84372 14266 84428
rect 14210 84292 14266 84348
rect 17100 84532 17156 84588
rect 17100 84452 17156 84508
rect 17100 84372 17156 84428
rect 17100 84292 17156 84348
rect 19990 84532 20046 84588
rect 19990 84452 20046 84508
rect 19990 84372 20046 84428
rect 19990 84292 20046 84348
rect 22880 84532 22936 84588
rect 22880 84452 22936 84508
rect 22880 84372 22936 84428
rect 22880 84292 22936 84348
rect 25770 84532 25826 84588
rect 25770 84452 25826 84508
rect 25770 84372 25826 84428
rect 25770 84292 25826 84348
rect 28660 84532 28716 84588
rect 28660 84452 28716 84508
rect 28660 84372 28716 84428
rect 28660 84292 28716 84348
rect 31550 84532 31606 84588
rect 31550 84452 31606 84508
rect 31550 84372 31606 84428
rect 31550 84292 31606 84348
rect 34440 84532 34496 84588
rect 34440 84452 34496 84508
rect 34440 84372 34496 84428
rect 34440 84292 34496 84348
rect 37330 84532 37386 84588
rect 37330 84452 37386 84508
rect 37330 84372 37386 84428
rect 37330 84292 37386 84348
rect 40220 84532 40276 84588
rect 40220 84452 40276 84508
rect 40220 84372 40276 84428
rect 40220 84292 40276 84348
rect 43110 84532 43166 84588
rect 43110 84452 43166 84508
rect 43110 84372 43166 84428
rect 43110 84292 43166 84348
rect 46000 84532 46056 84588
rect 46000 84452 46056 84508
rect 46000 84372 46056 84428
rect 46000 84292 46056 84348
rect 49008 84532 49064 84588
rect 49008 84452 49064 84508
rect 49008 84372 49064 84428
rect 49008 84292 49064 84348
rect 52237 84532 52293 84588
rect 52237 84452 52293 84508
rect 52237 84372 52293 84428
rect 52237 84292 52293 84348
rect 53638 84532 53694 84588
rect 53638 84452 53694 84508
rect 53638 84372 53694 84428
rect 53638 84292 53694 84348
rect 53806 84532 53862 84588
rect 53806 84452 53862 84508
rect 53806 84372 53862 84428
rect 53806 84292 53862 84348
rect 54550 84532 54606 84588
rect 54550 84452 54606 84508
rect 54550 84372 54606 84428
rect 54550 84292 54606 84348
rect 54940 84532 54996 84588
rect 54940 84452 54996 84508
rect 54940 84372 54996 84428
rect 54940 84292 54996 84348
rect 55656 84532 55712 84588
rect 55656 84452 55712 84508
rect 55656 84372 55712 84428
rect 55656 84292 55712 84348
rect 56234 84532 56290 84588
rect 56234 84452 56290 84508
rect 56234 84372 56290 84428
rect 56234 84292 56290 84348
rect 56679 84532 56735 84588
rect 56679 84452 56735 84508
rect 56679 84372 56735 84428
rect 56679 84292 56735 84348
rect 56983 84532 57039 84588
rect 56983 84452 57039 84508
rect 56983 84372 57039 84428
rect 56983 84292 57039 84348
rect 57825 84532 57881 84588
rect 57825 84452 57881 84508
rect 57825 84372 57881 84428
rect 57825 84292 57881 84348
rect 58465 84532 58521 84588
rect 58465 84452 58521 84508
rect 58465 84372 58521 84428
rect 58465 84292 58521 84348
rect 59048 84532 59104 84588
rect 59048 84452 59104 84508
rect 59048 84372 59104 84428
rect 59048 84292 59104 84348
rect 60326 84532 60382 84588
rect 60326 84452 60382 84508
rect 60326 84372 60382 84428
rect 60326 84292 60382 84348
rect 60484 84532 60540 84588
rect 60484 84452 60540 84508
rect 60484 84372 60540 84428
rect 60484 84292 60540 84348
rect 62528 84532 62584 84588
rect 62608 84532 62664 84588
rect 62528 84452 62584 84508
rect 62608 84452 62664 84508
rect 62528 84372 62584 84428
rect 62608 84372 62664 84428
rect 62528 84292 62584 84348
rect 62608 84292 62664 84348
rect 2184 82180 2240 82236
rect 2264 82180 2320 82236
rect 2184 82100 2240 82156
rect 2264 82100 2320 82156
rect 2184 82020 2240 82076
rect 2264 82020 2320 82076
rect 2184 81940 2240 81996
rect 2264 81940 2320 81996
rect 5393 82180 5449 82236
rect 5393 82100 5449 82156
rect 5393 82020 5449 82076
rect 5393 81940 5449 81996
rect 8283 82180 8339 82236
rect 8283 82100 8339 82156
rect 8283 82020 8339 82076
rect 8283 81940 8339 81996
rect 11173 82180 11229 82236
rect 11173 82100 11229 82156
rect 11173 82020 11229 82076
rect 11173 81940 11229 81996
rect 14063 82180 14119 82236
rect 14063 82100 14119 82156
rect 14063 82020 14119 82076
rect 14063 81940 14119 81996
rect 16953 82180 17009 82236
rect 16953 82100 17009 82156
rect 16953 82020 17009 82076
rect 16953 81940 17009 81996
rect 19843 82180 19899 82236
rect 19843 82100 19899 82156
rect 19843 82020 19899 82076
rect 19843 81940 19899 81996
rect 22733 82180 22789 82236
rect 22733 82100 22789 82156
rect 22733 82020 22789 82076
rect 22733 81940 22789 81996
rect 25623 82180 25679 82236
rect 25623 82100 25679 82156
rect 25623 82020 25679 82076
rect 25623 81940 25679 81996
rect 28513 82180 28569 82236
rect 28513 82100 28569 82156
rect 28513 82020 28569 82076
rect 28513 81940 28569 81996
rect 31403 82180 31459 82236
rect 31403 82100 31459 82156
rect 31403 82020 31459 82076
rect 31403 81940 31459 81996
rect 34293 82180 34349 82236
rect 34293 82100 34349 82156
rect 34293 82020 34349 82076
rect 34293 81940 34349 81996
rect 37183 82180 37239 82236
rect 37183 82100 37239 82156
rect 37183 82020 37239 82076
rect 37183 81940 37239 81996
rect 40073 82180 40129 82236
rect 40073 82100 40129 82156
rect 40073 82020 40129 82076
rect 40073 81940 40129 81996
rect 42963 82180 43019 82236
rect 42963 82100 43019 82156
rect 42963 82020 43019 82076
rect 42963 81940 43019 81996
rect 45853 82180 45909 82236
rect 45853 82100 45909 82156
rect 45853 82020 45909 82076
rect 45853 81940 45909 81996
rect 48800 82180 48856 82236
rect 48800 82100 48856 82156
rect 48800 82020 48856 82076
rect 48800 81940 48856 81996
rect 49662 82180 49718 82236
rect 49742 82180 49798 82236
rect 49662 82100 49718 82156
rect 49742 82100 49798 82156
rect 49662 82020 49718 82076
rect 49742 82020 49798 82076
rect 49662 81940 49718 81996
rect 49742 81940 49798 81996
rect 52956 82180 53012 82236
rect 52956 82100 53012 82156
rect 52956 82020 53012 82076
rect 52956 81940 53012 81996
rect 53114 82180 53170 82236
rect 53114 82100 53170 82156
rect 53114 82020 53170 82076
rect 53114 81940 53170 81996
rect 53470 82180 53526 82236
rect 53470 82100 53526 82156
rect 53470 82020 53526 82076
rect 53470 81940 53526 81996
rect 54788 82180 54844 82236
rect 54788 82100 54844 82156
rect 54788 82020 54844 82076
rect 54788 81940 54844 81996
rect 55381 82180 55437 82236
rect 55381 82100 55437 82156
rect 55381 82020 55437 82076
rect 55381 81940 55437 81996
rect 56527 82180 56583 82236
rect 56527 82100 56583 82156
rect 56527 82020 56583 82076
rect 56527 81940 56583 81996
rect 57963 82180 58019 82236
rect 58043 82180 58099 82236
rect 57963 82100 58019 82156
rect 58043 82100 58099 82156
rect 57963 82020 58019 82076
rect 58043 82020 58099 82076
rect 57963 81940 58019 81996
rect 58043 81940 58099 81996
rect 59206 82180 59262 82236
rect 59206 82100 59262 82156
rect 59206 82020 59262 82076
rect 59206 81940 59262 81996
rect 59364 82180 59420 82236
rect 59364 82100 59420 82156
rect 59364 82020 59420 82076
rect 59364 81940 59420 81996
rect 59672 82180 59728 82236
rect 59672 82100 59728 82156
rect 59672 82020 59728 82076
rect 59672 81940 59728 81996
rect 59818 82180 59874 82236
rect 59818 82100 59874 82156
rect 59818 82020 59874 82076
rect 59818 81940 59874 81996
rect 59954 82180 60010 82236
rect 60034 82180 60090 82236
rect 59954 82100 60010 82156
rect 60034 82100 60090 82156
rect 59954 82020 60010 82076
rect 60034 82020 60090 82076
rect 59954 81940 60010 81996
rect 60034 81940 60090 81996
rect 62326 82180 62382 82236
rect 62406 82180 62462 82236
rect 62326 82100 62382 82156
rect 62406 82100 62462 82156
rect 62326 82020 62382 82076
rect 62406 82020 62462 82076
rect 62326 81940 62382 81996
rect 62406 81940 62462 81996
rect 2044 74532 2100 74588
rect 2044 74452 2100 74508
rect 2044 74372 2100 74428
rect 2044 74292 2100 74348
rect 5540 74532 5596 74588
rect 5540 74452 5596 74508
rect 5540 74372 5596 74428
rect 5540 74292 5596 74348
rect 8430 74532 8486 74588
rect 8430 74452 8486 74508
rect 8430 74372 8486 74428
rect 8430 74292 8486 74348
rect 11320 74532 11376 74588
rect 11320 74452 11376 74508
rect 11320 74372 11376 74428
rect 11320 74292 11376 74348
rect 14210 74532 14266 74588
rect 14210 74452 14266 74508
rect 14210 74372 14266 74428
rect 14210 74292 14266 74348
rect 17100 74532 17156 74588
rect 17100 74452 17156 74508
rect 17100 74372 17156 74428
rect 17100 74292 17156 74348
rect 19990 74532 20046 74588
rect 19990 74452 20046 74508
rect 19990 74372 20046 74428
rect 19990 74292 20046 74348
rect 22880 74532 22936 74588
rect 22880 74452 22936 74508
rect 22880 74372 22936 74428
rect 22880 74292 22936 74348
rect 25770 74532 25826 74588
rect 25770 74452 25826 74508
rect 25770 74372 25826 74428
rect 25770 74292 25826 74348
rect 28660 74532 28716 74588
rect 28660 74452 28716 74508
rect 28660 74372 28716 74428
rect 28660 74292 28716 74348
rect 31550 74532 31606 74588
rect 31550 74452 31606 74508
rect 31550 74372 31606 74428
rect 31550 74292 31606 74348
rect 34440 74532 34496 74588
rect 34440 74452 34496 74508
rect 34440 74372 34496 74428
rect 34440 74292 34496 74348
rect 37330 74532 37386 74588
rect 37330 74452 37386 74508
rect 37330 74372 37386 74428
rect 37330 74292 37386 74348
rect 40220 74532 40276 74588
rect 40220 74452 40276 74508
rect 40220 74372 40276 74428
rect 40220 74292 40276 74348
rect 43110 74532 43166 74588
rect 43110 74452 43166 74508
rect 43110 74372 43166 74428
rect 43110 74292 43166 74348
rect 46000 74532 46056 74588
rect 46000 74452 46056 74508
rect 46000 74372 46056 74428
rect 46000 74292 46056 74348
rect 49008 74532 49064 74588
rect 49008 74452 49064 74508
rect 49008 74372 49064 74428
rect 49008 74292 49064 74348
rect 52237 74532 52293 74588
rect 52237 74452 52293 74508
rect 52237 74372 52293 74428
rect 52237 74292 52293 74348
rect 53638 74532 53694 74588
rect 53638 74452 53694 74508
rect 53638 74372 53694 74428
rect 53638 74292 53694 74348
rect 53806 74532 53862 74588
rect 53806 74452 53862 74508
rect 53806 74372 53862 74428
rect 53806 74292 53862 74348
rect 54550 74532 54606 74588
rect 54550 74452 54606 74508
rect 54550 74372 54606 74428
rect 54550 74292 54606 74348
rect 54940 74532 54996 74588
rect 54940 74452 54996 74508
rect 54940 74372 54996 74428
rect 54940 74292 54996 74348
rect 55656 74532 55712 74588
rect 55656 74452 55712 74508
rect 55656 74372 55712 74428
rect 55656 74292 55712 74348
rect 56234 74532 56290 74588
rect 56234 74452 56290 74508
rect 56234 74372 56290 74428
rect 56234 74292 56290 74348
rect 56679 74532 56735 74588
rect 56679 74452 56735 74508
rect 56679 74372 56735 74428
rect 56679 74292 56735 74348
rect 56983 74532 57039 74588
rect 56983 74452 57039 74508
rect 56983 74372 57039 74428
rect 56983 74292 57039 74348
rect 57825 74532 57881 74588
rect 57825 74452 57881 74508
rect 57825 74372 57881 74428
rect 57825 74292 57881 74348
rect 58465 74532 58521 74588
rect 58465 74452 58521 74508
rect 58465 74372 58521 74428
rect 58465 74292 58521 74348
rect 59048 74532 59104 74588
rect 59048 74452 59104 74508
rect 59048 74372 59104 74428
rect 59048 74292 59104 74348
rect 60326 74532 60382 74588
rect 60326 74452 60382 74508
rect 60326 74372 60382 74428
rect 60326 74292 60382 74348
rect 60484 74532 60540 74588
rect 60484 74452 60540 74508
rect 60484 74372 60540 74428
rect 60484 74292 60540 74348
rect 62528 74532 62584 74588
rect 62608 74532 62664 74588
rect 62528 74452 62584 74508
rect 62608 74452 62664 74508
rect 62528 74372 62584 74428
rect 62608 74372 62664 74428
rect 62528 74292 62584 74348
rect 62608 74292 62664 74348
rect 2184 72180 2240 72236
rect 2264 72180 2320 72236
rect 2184 72100 2240 72156
rect 2264 72100 2320 72156
rect 2184 72020 2240 72076
rect 2264 72020 2320 72076
rect 2184 71940 2240 71996
rect 2264 71940 2320 71996
rect 5393 72180 5449 72236
rect 5393 72100 5449 72156
rect 5393 72020 5449 72076
rect 5393 71940 5449 71996
rect 8283 72180 8339 72236
rect 8283 72100 8339 72156
rect 8283 72020 8339 72076
rect 8283 71940 8339 71996
rect 11173 72180 11229 72236
rect 11173 72100 11229 72156
rect 11173 72020 11229 72076
rect 11173 71940 11229 71996
rect 14063 72180 14119 72236
rect 14063 72100 14119 72156
rect 14063 72020 14119 72076
rect 14063 71940 14119 71996
rect 16953 72180 17009 72236
rect 16953 72100 17009 72156
rect 16953 72020 17009 72076
rect 16953 71940 17009 71996
rect 19843 72180 19899 72236
rect 19843 72100 19899 72156
rect 19843 72020 19899 72076
rect 19843 71940 19899 71996
rect 22733 72180 22789 72236
rect 22733 72100 22789 72156
rect 22733 72020 22789 72076
rect 22733 71940 22789 71996
rect 25623 72180 25679 72236
rect 25623 72100 25679 72156
rect 25623 72020 25679 72076
rect 25623 71940 25679 71996
rect 28513 72180 28569 72236
rect 28513 72100 28569 72156
rect 28513 72020 28569 72076
rect 28513 71940 28569 71996
rect 31403 72180 31459 72236
rect 31403 72100 31459 72156
rect 31403 72020 31459 72076
rect 31403 71940 31459 71996
rect 34293 72180 34349 72236
rect 34293 72100 34349 72156
rect 34293 72020 34349 72076
rect 34293 71940 34349 71996
rect 37183 72180 37239 72236
rect 37183 72100 37239 72156
rect 37183 72020 37239 72076
rect 37183 71940 37239 71996
rect 40073 72180 40129 72236
rect 40073 72100 40129 72156
rect 40073 72020 40129 72076
rect 40073 71940 40129 71996
rect 42963 72180 43019 72236
rect 42963 72100 43019 72156
rect 42963 72020 43019 72076
rect 42963 71940 43019 71996
rect 45853 72180 45909 72236
rect 45853 72100 45909 72156
rect 45853 72020 45909 72076
rect 45853 71940 45909 71996
rect 48800 72180 48856 72236
rect 48800 72100 48856 72156
rect 48800 72020 48856 72076
rect 48800 71940 48856 71996
rect 49662 72180 49718 72236
rect 49742 72180 49798 72236
rect 49662 72100 49718 72156
rect 49742 72100 49798 72156
rect 49662 72020 49718 72076
rect 49742 72020 49798 72076
rect 49662 71940 49718 71996
rect 49742 71940 49798 71996
rect 52956 72180 53012 72236
rect 52956 72100 53012 72156
rect 52956 72020 53012 72076
rect 52956 71940 53012 71996
rect 53114 72180 53170 72236
rect 53114 72100 53170 72156
rect 53114 72020 53170 72076
rect 53114 71940 53170 71996
rect 53470 72180 53526 72236
rect 53470 72100 53526 72156
rect 53470 72020 53526 72076
rect 53470 71940 53526 71996
rect 54788 72180 54844 72236
rect 54788 72100 54844 72156
rect 54788 72020 54844 72076
rect 54788 71940 54844 71996
rect 55381 72180 55437 72236
rect 55381 72100 55437 72156
rect 55381 72020 55437 72076
rect 55381 71940 55437 71996
rect 56527 72180 56583 72236
rect 56527 72100 56583 72156
rect 56527 72020 56583 72076
rect 56527 71940 56583 71996
rect 57963 72180 58019 72236
rect 58043 72180 58099 72236
rect 57963 72100 58019 72156
rect 58043 72100 58099 72156
rect 57963 72020 58019 72076
rect 58043 72020 58099 72076
rect 57963 71940 58019 71996
rect 58043 71940 58099 71996
rect 59206 72180 59262 72236
rect 59206 72100 59262 72156
rect 59206 72020 59262 72076
rect 59206 71940 59262 71996
rect 59364 72180 59420 72236
rect 59364 72100 59420 72156
rect 59364 72020 59420 72076
rect 59364 71940 59420 71996
rect 59672 72180 59728 72236
rect 59672 72100 59728 72156
rect 59672 72020 59728 72076
rect 59672 71940 59728 71996
rect 59818 72180 59874 72236
rect 59818 72100 59874 72156
rect 59818 72020 59874 72076
rect 59818 71940 59874 71996
rect 59954 72180 60010 72236
rect 60034 72180 60090 72236
rect 59954 72100 60010 72156
rect 60034 72100 60090 72156
rect 59954 72020 60010 72076
rect 60034 72020 60090 72076
rect 59954 71940 60010 71996
rect 60034 71940 60090 71996
rect 62326 72180 62382 72236
rect 62406 72180 62462 72236
rect 62326 72100 62382 72156
rect 62406 72100 62462 72156
rect 62326 72020 62382 72076
rect 62406 72020 62462 72076
rect 62326 71940 62382 71996
rect 62406 71940 62462 71996
rect 2044 64532 2100 64588
rect 2044 64452 2100 64508
rect 2044 64372 2100 64428
rect 2044 64292 2100 64348
rect 5540 64532 5596 64588
rect 5540 64452 5596 64508
rect 5540 64372 5596 64428
rect 5540 64292 5596 64348
rect 8430 64532 8486 64588
rect 8430 64452 8486 64508
rect 8430 64372 8486 64428
rect 8430 64292 8486 64348
rect 11320 64532 11376 64588
rect 11320 64452 11376 64508
rect 11320 64372 11376 64428
rect 11320 64292 11376 64348
rect 14210 64532 14266 64588
rect 14210 64452 14266 64508
rect 14210 64372 14266 64428
rect 14210 64292 14266 64348
rect 17100 64532 17156 64588
rect 17100 64452 17156 64508
rect 17100 64372 17156 64428
rect 17100 64292 17156 64348
rect 19990 64532 20046 64588
rect 19990 64452 20046 64508
rect 19990 64372 20046 64428
rect 19990 64292 20046 64348
rect 22880 64532 22936 64588
rect 22880 64452 22936 64508
rect 22880 64372 22936 64428
rect 22880 64292 22936 64348
rect 25770 64532 25826 64588
rect 25770 64452 25826 64508
rect 25770 64372 25826 64428
rect 25770 64292 25826 64348
rect 28660 64532 28716 64588
rect 28660 64452 28716 64508
rect 28660 64372 28716 64428
rect 28660 64292 28716 64348
rect 31550 64532 31606 64588
rect 31550 64452 31606 64508
rect 31550 64372 31606 64428
rect 31550 64292 31606 64348
rect 34440 64532 34496 64588
rect 34440 64452 34496 64508
rect 34440 64372 34496 64428
rect 34440 64292 34496 64348
rect 37330 64532 37386 64588
rect 37330 64452 37386 64508
rect 37330 64372 37386 64428
rect 37330 64292 37386 64348
rect 40220 64532 40276 64588
rect 40220 64452 40276 64508
rect 40220 64372 40276 64428
rect 40220 64292 40276 64348
rect 43110 64532 43166 64588
rect 43110 64452 43166 64508
rect 43110 64372 43166 64428
rect 43110 64292 43166 64348
rect 46000 64532 46056 64588
rect 46000 64452 46056 64508
rect 46000 64372 46056 64428
rect 46000 64292 46056 64348
rect 49008 64532 49064 64588
rect 49008 64452 49064 64508
rect 49008 64372 49064 64428
rect 49008 64292 49064 64348
rect 52237 64532 52293 64588
rect 52237 64452 52293 64508
rect 52237 64372 52293 64428
rect 52237 64292 52293 64348
rect 53638 64532 53694 64588
rect 53638 64452 53694 64508
rect 53638 64372 53694 64428
rect 53638 64292 53694 64348
rect 53806 64532 53862 64588
rect 53806 64452 53862 64508
rect 53806 64372 53862 64428
rect 53806 64292 53862 64348
rect 54550 64532 54606 64588
rect 54550 64452 54606 64508
rect 54550 64372 54606 64428
rect 54550 64292 54606 64348
rect 54940 64532 54996 64588
rect 54940 64452 54996 64508
rect 54940 64372 54996 64428
rect 54940 64292 54996 64348
rect 55656 64532 55712 64588
rect 55656 64452 55712 64508
rect 55656 64372 55712 64428
rect 55656 64292 55712 64348
rect 56234 64532 56290 64588
rect 56234 64452 56290 64508
rect 56234 64372 56290 64428
rect 56234 64292 56290 64348
rect 56679 64532 56735 64588
rect 56679 64452 56735 64508
rect 56679 64372 56735 64428
rect 56679 64292 56735 64348
rect 56983 64532 57039 64588
rect 56983 64452 57039 64508
rect 56983 64372 57039 64428
rect 56983 64292 57039 64348
rect 57825 64532 57881 64588
rect 57825 64452 57881 64508
rect 57825 64372 57881 64428
rect 57825 64292 57881 64348
rect 58465 64532 58521 64588
rect 58465 64452 58521 64508
rect 58465 64372 58521 64428
rect 58465 64292 58521 64348
rect 59048 64532 59104 64588
rect 59048 64452 59104 64508
rect 59048 64372 59104 64428
rect 59048 64292 59104 64348
rect 60326 64532 60382 64588
rect 60326 64452 60382 64508
rect 60326 64372 60382 64428
rect 60326 64292 60382 64348
rect 60484 64532 60540 64588
rect 60484 64452 60540 64508
rect 60484 64372 60540 64428
rect 60484 64292 60540 64348
rect 62528 64532 62584 64588
rect 62608 64532 62664 64588
rect 62528 64452 62584 64508
rect 62608 64452 62664 64508
rect 62528 64372 62584 64428
rect 62608 64372 62664 64428
rect 62528 64292 62584 64348
rect 62608 64292 62664 64348
rect 2184 62180 2240 62236
rect 2264 62180 2320 62236
rect 2184 62100 2240 62156
rect 2264 62100 2320 62156
rect 2184 62020 2240 62076
rect 2264 62020 2320 62076
rect 2184 61940 2240 61996
rect 2264 61940 2320 61996
rect 5393 62180 5449 62236
rect 5393 62100 5449 62156
rect 5393 62020 5449 62076
rect 5393 61940 5449 61996
rect 8283 62180 8339 62236
rect 8283 62100 8339 62156
rect 8283 62020 8339 62076
rect 8283 61940 8339 61996
rect 11173 62180 11229 62236
rect 11173 62100 11229 62156
rect 11173 62020 11229 62076
rect 11173 61940 11229 61996
rect 14063 62180 14119 62236
rect 14063 62100 14119 62156
rect 14063 62020 14119 62076
rect 14063 61940 14119 61996
rect 16953 62180 17009 62236
rect 16953 62100 17009 62156
rect 16953 62020 17009 62076
rect 16953 61940 17009 61996
rect 19843 62180 19899 62236
rect 19843 62100 19899 62156
rect 19843 62020 19899 62076
rect 19843 61940 19899 61996
rect 22733 62180 22789 62236
rect 22733 62100 22789 62156
rect 22733 62020 22789 62076
rect 22733 61940 22789 61996
rect 25623 62180 25679 62236
rect 25623 62100 25679 62156
rect 25623 62020 25679 62076
rect 25623 61940 25679 61996
rect 28513 62180 28569 62236
rect 28513 62100 28569 62156
rect 28513 62020 28569 62076
rect 28513 61940 28569 61996
rect 31403 62180 31459 62236
rect 31403 62100 31459 62156
rect 31403 62020 31459 62076
rect 31403 61940 31459 61996
rect 34293 62180 34349 62236
rect 34293 62100 34349 62156
rect 34293 62020 34349 62076
rect 34293 61940 34349 61996
rect 37183 62180 37239 62236
rect 37183 62100 37239 62156
rect 37183 62020 37239 62076
rect 37183 61940 37239 61996
rect 40073 62180 40129 62236
rect 40073 62100 40129 62156
rect 40073 62020 40129 62076
rect 40073 61940 40129 61996
rect 42963 62180 43019 62236
rect 42963 62100 43019 62156
rect 42963 62020 43019 62076
rect 42963 61940 43019 61996
rect 45853 62180 45909 62236
rect 45853 62100 45909 62156
rect 45853 62020 45909 62076
rect 45853 61940 45909 61996
rect 48800 62180 48856 62236
rect 48800 62100 48856 62156
rect 48800 62020 48856 62076
rect 48800 61940 48856 61996
rect 49662 62180 49718 62236
rect 49742 62180 49798 62236
rect 49662 62100 49718 62156
rect 49742 62100 49798 62156
rect 49662 62020 49718 62076
rect 49742 62020 49798 62076
rect 49662 61940 49718 61996
rect 49742 61940 49798 61996
rect 52956 62180 53012 62236
rect 52956 62100 53012 62156
rect 52956 62020 53012 62076
rect 52956 61940 53012 61996
rect 53114 62180 53170 62236
rect 53114 62100 53170 62156
rect 53114 62020 53170 62076
rect 53114 61940 53170 61996
rect 53470 62180 53526 62236
rect 53470 62100 53526 62156
rect 53470 62020 53526 62076
rect 53470 61940 53526 61996
rect 54788 62180 54844 62236
rect 54788 62100 54844 62156
rect 54788 62020 54844 62076
rect 54788 61940 54844 61996
rect 55381 62180 55437 62236
rect 55381 62100 55437 62156
rect 55381 62020 55437 62076
rect 55381 61940 55437 61996
rect 56527 62180 56583 62236
rect 56527 62100 56583 62156
rect 56527 62020 56583 62076
rect 56527 61940 56583 61996
rect 57963 62180 58019 62236
rect 58043 62180 58099 62236
rect 57963 62100 58019 62156
rect 58043 62100 58099 62156
rect 57963 62020 58019 62076
rect 58043 62020 58099 62076
rect 57963 61940 58019 61996
rect 58043 61940 58099 61996
rect 59206 62180 59262 62236
rect 59206 62100 59262 62156
rect 59206 62020 59262 62076
rect 59206 61940 59262 61996
rect 59364 62180 59420 62236
rect 59364 62100 59420 62156
rect 59364 62020 59420 62076
rect 59364 61940 59420 61996
rect 59672 62180 59728 62236
rect 59672 62100 59728 62156
rect 59672 62020 59728 62076
rect 59672 61940 59728 61996
rect 59818 62180 59874 62236
rect 59818 62100 59874 62156
rect 59818 62020 59874 62076
rect 59818 61940 59874 61996
rect 59954 62180 60010 62236
rect 60034 62180 60090 62236
rect 59954 62100 60010 62156
rect 60034 62100 60090 62156
rect 59954 62020 60010 62076
rect 60034 62020 60090 62076
rect 59954 61940 60010 61996
rect 60034 61940 60090 61996
rect 62326 62180 62382 62236
rect 62406 62180 62462 62236
rect 62326 62100 62382 62156
rect 62406 62100 62462 62156
rect 62326 62020 62382 62076
rect 62406 62020 62462 62076
rect 62326 61940 62382 61996
rect 62406 61940 62462 61996
rect 2044 54532 2100 54588
rect 2044 54452 2100 54508
rect 2044 54372 2100 54428
rect 2044 54292 2100 54348
rect 5540 54532 5596 54588
rect 5540 54452 5596 54508
rect 5540 54372 5596 54428
rect 5540 54292 5596 54348
rect 8430 54532 8486 54588
rect 8430 54452 8486 54508
rect 8430 54372 8486 54428
rect 8430 54292 8486 54348
rect 11320 54532 11376 54588
rect 11320 54452 11376 54508
rect 11320 54372 11376 54428
rect 11320 54292 11376 54348
rect 14210 54532 14266 54588
rect 14210 54452 14266 54508
rect 14210 54372 14266 54428
rect 14210 54292 14266 54348
rect 17100 54532 17156 54588
rect 17100 54452 17156 54508
rect 17100 54372 17156 54428
rect 17100 54292 17156 54348
rect 19990 54532 20046 54588
rect 19990 54452 20046 54508
rect 19990 54372 20046 54428
rect 19990 54292 20046 54348
rect 22880 54532 22936 54588
rect 22880 54452 22936 54508
rect 22880 54372 22936 54428
rect 22880 54292 22936 54348
rect 25770 54532 25826 54588
rect 25770 54452 25826 54508
rect 25770 54372 25826 54428
rect 25770 54292 25826 54348
rect 28660 54532 28716 54588
rect 28660 54452 28716 54508
rect 28660 54372 28716 54428
rect 28660 54292 28716 54348
rect 31550 54532 31606 54588
rect 31550 54452 31606 54508
rect 31550 54372 31606 54428
rect 31550 54292 31606 54348
rect 34440 54532 34496 54588
rect 34440 54452 34496 54508
rect 34440 54372 34496 54428
rect 34440 54292 34496 54348
rect 37330 54532 37386 54588
rect 37330 54452 37386 54508
rect 37330 54372 37386 54428
rect 37330 54292 37386 54348
rect 40220 54532 40276 54588
rect 40220 54452 40276 54508
rect 40220 54372 40276 54428
rect 40220 54292 40276 54348
rect 43110 54532 43166 54588
rect 43110 54452 43166 54508
rect 43110 54372 43166 54428
rect 43110 54292 43166 54348
rect 46000 54532 46056 54588
rect 46000 54452 46056 54508
rect 46000 54372 46056 54428
rect 46000 54292 46056 54348
rect 49008 54532 49064 54588
rect 49008 54452 49064 54508
rect 49008 54372 49064 54428
rect 49008 54292 49064 54348
rect 52237 54532 52293 54588
rect 52237 54452 52293 54508
rect 52237 54372 52293 54428
rect 52237 54292 52293 54348
rect 53638 54532 53694 54588
rect 53638 54452 53694 54508
rect 53638 54372 53694 54428
rect 53638 54292 53694 54348
rect 53806 54532 53862 54588
rect 53806 54452 53862 54508
rect 53806 54372 53862 54428
rect 53806 54292 53862 54348
rect 54550 54532 54606 54588
rect 54550 54452 54606 54508
rect 54550 54372 54606 54428
rect 54550 54292 54606 54348
rect 54940 54532 54996 54588
rect 54940 54452 54996 54508
rect 54940 54372 54996 54428
rect 54940 54292 54996 54348
rect 55656 54532 55712 54588
rect 55656 54452 55712 54508
rect 55656 54372 55712 54428
rect 55656 54292 55712 54348
rect 56234 54532 56290 54588
rect 56234 54452 56290 54508
rect 56234 54372 56290 54428
rect 56234 54292 56290 54348
rect 56679 54532 56735 54588
rect 56679 54452 56735 54508
rect 56679 54372 56735 54428
rect 56679 54292 56735 54348
rect 56983 54532 57039 54588
rect 56983 54452 57039 54508
rect 56983 54372 57039 54428
rect 56983 54292 57039 54348
rect 57825 54532 57881 54588
rect 57825 54452 57881 54508
rect 57825 54372 57881 54428
rect 57825 54292 57881 54348
rect 58465 54532 58521 54588
rect 58465 54452 58521 54508
rect 58465 54372 58521 54428
rect 58465 54292 58521 54348
rect 59048 54532 59104 54588
rect 59048 54452 59104 54508
rect 59048 54372 59104 54428
rect 59048 54292 59104 54348
rect 60326 54532 60382 54588
rect 60326 54452 60382 54508
rect 60326 54372 60382 54428
rect 60326 54292 60382 54348
rect 60484 54532 60540 54588
rect 60484 54452 60540 54508
rect 60484 54372 60540 54428
rect 60484 54292 60540 54348
rect 62528 54532 62584 54588
rect 62608 54532 62664 54588
rect 62528 54452 62584 54508
rect 62608 54452 62664 54508
rect 62528 54372 62584 54428
rect 62608 54372 62664 54428
rect 62528 54292 62584 54348
rect 62608 54292 62664 54348
rect 2184 52180 2240 52236
rect 2264 52180 2320 52236
rect 2184 52100 2240 52156
rect 2264 52100 2320 52156
rect 2184 52020 2240 52076
rect 2264 52020 2320 52076
rect 2184 51940 2240 51996
rect 2264 51940 2320 51996
rect 5393 52180 5449 52236
rect 5393 52100 5449 52156
rect 5393 52020 5449 52076
rect 5393 51940 5449 51996
rect 8283 52180 8339 52236
rect 8283 52100 8339 52156
rect 8283 52020 8339 52076
rect 8283 51940 8339 51996
rect 11173 52180 11229 52236
rect 11173 52100 11229 52156
rect 11173 52020 11229 52076
rect 11173 51940 11229 51996
rect 14063 52180 14119 52236
rect 14063 52100 14119 52156
rect 14063 52020 14119 52076
rect 14063 51940 14119 51996
rect 16953 52180 17009 52236
rect 16953 52100 17009 52156
rect 16953 52020 17009 52076
rect 16953 51940 17009 51996
rect 19843 52180 19899 52236
rect 19843 52100 19899 52156
rect 19843 52020 19899 52076
rect 19843 51940 19899 51996
rect 22733 52180 22789 52236
rect 22733 52100 22789 52156
rect 22733 52020 22789 52076
rect 22733 51940 22789 51996
rect 25623 52180 25679 52236
rect 25623 52100 25679 52156
rect 25623 52020 25679 52076
rect 25623 51940 25679 51996
rect 28513 52180 28569 52236
rect 28513 52100 28569 52156
rect 28513 52020 28569 52076
rect 28513 51940 28569 51996
rect 31403 52180 31459 52236
rect 31403 52100 31459 52156
rect 31403 52020 31459 52076
rect 31403 51940 31459 51996
rect 34293 52180 34349 52236
rect 34293 52100 34349 52156
rect 34293 52020 34349 52076
rect 34293 51940 34349 51996
rect 37183 52180 37239 52236
rect 37183 52100 37239 52156
rect 37183 52020 37239 52076
rect 37183 51940 37239 51996
rect 40073 52180 40129 52236
rect 40073 52100 40129 52156
rect 40073 52020 40129 52076
rect 40073 51940 40129 51996
rect 42963 52180 43019 52236
rect 42963 52100 43019 52156
rect 42963 52020 43019 52076
rect 42963 51940 43019 51996
rect 45853 52180 45909 52236
rect 45853 52100 45909 52156
rect 45853 52020 45909 52076
rect 45853 51940 45909 51996
rect 48800 52180 48856 52236
rect 48800 52100 48856 52156
rect 48800 52020 48856 52076
rect 48800 51940 48856 51996
rect 49662 52180 49718 52236
rect 49742 52180 49798 52236
rect 49662 52100 49718 52156
rect 49742 52100 49798 52156
rect 49662 52020 49718 52076
rect 49742 52020 49798 52076
rect 49662 51940 49718 51996
rect 49742 51940 49798 51996
rect 52956 52180 53012 52236
rect 52956 52100 53012 52156
rect 52956 52020 53012 52076
rect 52956 51940 53012 51996
rect 53114 52180 53170 52236
rect 53114 52100 53170 52156
rect 53114 52020 53170 52076
rect 53114 51940 53170 51996
rect 53470 52180 53526 52236
rect 53470 52100 53526 52156
rect 53470 52020 53526 52076
rect 53470 51940 53526 51996
rect 54788 52180 54844 52236
rect 54788 52100 54844 52156
rect 54788 52020 54844 52076
rect 54788 51940 54844 51996
rect 55381 52180 55437 52236
rect 55381 52100 55437 52156
rect 55381 52020 55437 52076
rect 55381 51940 55437 51996
rect 56527 52180 56583 52236
rect 56527 52100 56583 52156
rect 56527 52020 56583 52076
rect 56527 51940 56583 51996
rect 57963 52180 58019 52236
rect 58043 52180 58099 52236
rect 57963 52100 58019 52156
rect 58043 52100 58099 52156
rect 57963 52020 58019 52076
rect 58043 52020 58099 52076
rect 57963 51940 58019 51996
rect 58043 51940 58099 51996
rect 59206 52180 59262 52236
rect 59206 52100 59262 52156
rect 59206 52020 59262 52076
rect 59206 51940 59262 51996
rect 59364 52180 59420 52236
rect 59364 52100 59420 52156
rect 59364 52020 59420 52076
rect 59364 51940 59420 51996
rect 59672 52180 59728 52236
rect 59672 52100 59728 52156
rect 59672 52020 59728 52076
rect 59672 51940 59728 51996
rect 59818 52180 59874 52236
rect 59818 52100 59874 52156
rect 59818 52020 59874 52076
rect 59818 51940 59874 51996
rect 59954 52180 60010 52236
rect 60034 52180 60090 52236
rect 59954 52100 60010 52156
rect 60034 52100 60090 52156
rect 59954 52020 60010 52076
rect 60034 52020 60090 52076
rect 59954 51940 60010 51996
rect 60034 51940 60090 51996
rect 62326 52180 62382 52236
rect 62406 52180 62462 52236
rect 62326 52100 62382 52156
rect 62406 52100 62462 52156
rect 62326 52020 62382 52076
rect 62406 52020 62462 52076
rect 62326 51940 62382 51996
rect 62406 51940 62462 51996
rect 2044 44532 2100 44588
rect 2044 44452 2100 44508
rect 2044 44372 2100 44428
rect 2044 44292 2100 44348
rect 5540 44532 5596 44588
rect 5540 44452 5596 44508
rect 5540 44372 5596 44428
rect 5540 44292 5596 44348
rect 8430 44532 8486 44588
rect 8430 44452 8486 44508
rect 8430 44372 8486 44428
rect 8430 44292 8486 44348
rect 11320 44532 11376 44588
rect 11320 44452 11376 44508
rect 11320 44372 11376 44428
rect 11320 44292 11376 44348
rect 14210 44532 14266 44588
rect 14210 44452 14266 44508
rect 14210 44372 14266 44428
rect 14210 44292 14266 44348
rect 17100 44532 17156 44588
rect 17100 44452 17156 44508
rect 17100 44372 17156 44428
rect 17100 44292 17156 44348
rect 19990 44532 20046 44588
rect 19990 44452 20046 44508
rect 19990 44372 20046 44428
rect 19990 44292 20046 44348
rect 22880 44532 22936 44588
rect 22880 44452 22936 44508
rect 22880 44372 22936 44428
rect 22880 44292 22936 44348
rect 25770 44532 25826 44588
rect 25770 44452 25826 44508
rect 25770 44372 25826 44428
rect 25770 44292 25826 44348
rect 28660 44532 28716 44588
rect 28660 44452 28716 44508
rect 28660 44372 28716 44428
rect 28660 44292 28716 44348
rect 31550 44532 31606 44588
rect 31550 44452 31606 44508
rect 31550 44372 31606 44428
rect 31550 44292 31606 44348
rect 34440 44532 34496 44588
rect 34440 44452 34496 44508
rect 34440 44372 34496 44428
rect 34440 44292 34496 44348
rect 37330 44532 37386 44588
rect 37330 44452 37386 44508
rect 37330 44372 37386 44428
rect 37330 44292 37386 44348
rect 40220 44532 40276 44588
rect 40220 44452 40276 44508
rect 40220 44372 40276 44428
rect 40220 44292 40276 44348
rect 43110 44532 43166 44588
rect 43110 44452 43166 44508
rect 43110 44372 43166 44428
rect 43110 44292 43166 44348
rect 46000 44532 46056 44588
rect 46000 44452 46056 44508
rect 46000 44372 46056 44428
rect 46000 44292 46056 44348
rect 52237 44532 52293 44588
rect 52237 44452 52293 44508
rect 52237 44372 52293 44428
rect 52237 44292 52293 44348
rect 53638 44532 53694 44588
rect 53638 44452 53694 44508
rect 53638 44372 53694 44428
rect 53638 44292 53694 44348
rect 54550 44532 54606 44588
rect 54550 44452 54606 44508
rect 54550 44372 54606 44428
rect 54550 44292 54606 44348
rect 54940 44532 54996 44588
rect 54940 44452 54996 44508
rect 54940 44372 54996 44428
rect 54940 44292 54996 44348
rect 55656 44532 55712 44588
rect 55656 44452 55712 44508
rect 55656 44372 55712 44428
rect 55656 44292 55712 44348
rect 56234 44532 56290 44588
rect 56234 44452 56290 44508
rect 56234 44372 56290 44428
rect 56234 44292 56290 44348
rect 56679 44532 56735 44588
rect 56679 44452 56735 44508
rect 56679 44372 56735 44428
rect 56679 44292 56735 44348
rect 56983 44532 57039 44588
rect 56983 44452 57039 44508
rect 56983 44372 57039 44428
rect 56983 44292 57039 44348
rect 57825 44532 57881 44588
rect 57825 44452 57881 44508
rect 57825 44372 57881 44428
rect 57825 44292 57881 44348
rect 58349 44532 58405 44588
rect 58349 44452 58405 44508
rect 58349 44372 58405 44428
rect 58349 44292 58405 44348
rect 59048 44532 59104 44588
rect 59048 44452 59104 44508
rect 59048 44372 59104 44428
rect 59048 44292 59104 44348
rect 60326 44532 60382 44588
rect 60326 44452 60382 44508
rect 60326 44372 60382 44428
rect 60326 44292 60382 44348
rect 60484 44532 60540 44588
rect 60484 44452 60540 44508
rect 60484 44372 60540 44428
rect 60484 44292 60540 44348
rect 62528 44532 62584 44588
rect 62608 44532 62664 44588
rect 62528 44452 62584 44508
rect 62608 44452 62664 44508
rect 62528 44372 62584 44428
rect 62608 44372 62664 44428
rect 62528 44292 62584 44348
rect 62608 44292 62664 44348
rect 2184 42180 2240 42236
rect 2264 42180 2320 42236
rect 2184 42100 2240 42156
rect 2264 42100 2320 42156
rect 2184 42020 2240 42076
rect 2264 42020 2320 42076
rect 2184 41940 2240 41996
rect 2264 41940 2320 41996
rect 5393 42180 5449 42236
rect 5393 42100 5449 42156
rect 5393 42020 5449 42076
rect 5393 41940 5449 41996
rect 8283 42180 8339 42236
rect 8283 42100 8339 42156
rect 8283 42020 8339 42076
rect 8283 41940 8339 41996
rect 11173 42180 11229 42236
rect 11173 42100 11229 42156
rect 11173 42020 11229 42076
rect 11173 41940 11229 41996
rect 14063 42180 14119 42236
rect 14063 42100 14119 42156
rect 14063 42020 14119 42076
rect 14063 41940 14119 41996
rect 16953 42180 17009 42236
rect 16953 42100 17009 42156
rect 16953 42020 17009 42076
rect 16953 41940 17009 41996
rect 19843 42180 19899 42236
rect 19843 42100 19899 42156
rect 19843 42020 19899 42076
rect 19843 41940 19899 41996
rect 22733 42180 22789 42236
rect 22733 42100 22789 42156
rect 22733 42020 22789 42076
rect 22733 41940 22789 41996
rect 25623 42180 25679 42236
rect 25623 42100 25679 42156
rect 25623 42020 25679 42076
rect 25623 41940 25679 41996
rect 28513 42180 28569 42236
rect 28513 42100 28569 42156
rect 28513 42020 28569 42076
rect 28513 41940 28569 41996
rect 31403 42180 31459 42236
rect 31403 42100 31459 42156
rect 31403 42020 31459 42076
rect 31403 41940 31459 41996
rect 34293 42180 34349 42236
rect 34293 42100 34349 42156
rect 34293 42020 34349 42076
rect 34293 41940 34349 41996
rect 37183 42180 37239 42236
rect 37183 42100 37239 42156
rect 37183 42020 37239 42076
rect 37183 41940 37239 41996
rect 40073 42180 40129 42236
rect 40073 42100 40129 42156
rect 40073 42020 40129 42076
rect 40073 41940 40129 41996
rect 42963 42180 43019 42236
rect 42963 42100 43019 42156
rect 42963 42020 43019 42076
rect 42963 41940 43019 41996
rect 45853 42180 45909 42236
rect 45853 42100 45909 42156
rect 45853 42020 45909 42076
rect 45853 41940 45909 41996
rect 48800 42180 48856 42236
rect 48800 42100 48856 42156
rect 48800 42020 48856 42076
rect 48800 41940 48856 41996
rect 49662 42180 49718 42236
rect 49742 42180 49798 42236
rect 49662 42100 49718 42156
rect 49742 42100 49798 42156
rect 49662 42020 49718 42076
rect 49742 42020 49798 42076
rect 49662 41940 49718 41996
rect 49742 41940 49798 41996
rect 52956 42180 53012 42236
rect 52956 42100 53012 42156
rect 52956 42020 53012 42076
rect 52956 41940 53012 41996
rect 53114 42180 53170 42236
rect 53114 42100 53170 42156
rect 53114 42020 53170 42076
rect 53114 41940 53170 41996
rect 53470 42180 53526 42236
rect 53470 42100 53526 42156
rect 53470 42020 53526 42076
rect 53470 41940 53526 41996
rect 54788 42180 54844 42236
rect 54788 42100 54844 42156
rect 54788 42020 54844 42076
rect 54788 41940 54844 41996
rect 55381 42180 55437 42236
rect 55381 42100 55437 42156
rect 55381 42020 55437 42076
rect 55381 41940 55437 41996
rect 56527 42180 56583 42236
rect 56527 42100 56583 42156
rect 56527 42020 56583 42076
rect 56527 41940 56583 41996
rect 57963 42180 58019 42236
rect 58043 42180 58099 42236
rect 57963 42100 58019 42156
rect 58043 42100 58099 42156
rect 57963 42020 58019 42076
rect 58043 42020 58099 42076
rect 57963 41940 58019 41996
rect 58043 41940 58099 41996
rect 59206 42180 59262 42236
rect 59206 42100 59262 42156
rect 59206 42020 59262 42076
rect 59206 41940 59262 41996
rect 59364 42180 59420 42236
rect 59364 42100 59420 42156
rect 59364 42020 59420 42076
rect 59364 41940 59420 41996
rect 59672 42180 59728 42236
rect 59672 42100 59728 42156
rect 59672 42020 59728 42076
rect 59672 41940 59728 41996
rect 59818 42180 59874 42236
rect 59818 42100 59874 42156
rect 59818 42020 59874 42076
rect 59818 41940 59874 41996
rect 59954 42180 60010 42236
rect 60034 42180 60090 42236
rect 59954 42100 60010 42156
rect 60034 42100 60090 42156
rect 59954 42020 60010 42076
rect 60034 42020 60090 42076
rect 59954 41940 60010 41996
rect 60034 41940 60090 41996
rect 62326 42180 62382 42236
rect 62406 42180 62462 42236
rect 62326 42100 62382 42156
rect 62406 42100 62462 42156
rect 62326 42020 62382 42076
rect 62406 42020 62462 42076
rect 62326 41940 62382 41996
rect 62406 41940 62462 41996
rect 2044 34532 2100 34588
rect 2044 34452 2100 34508
rect 2044 34372 2100 34428
rect 2044 34292 2100 34348
rect 5540 34532 5596 34588
rect 5540 34452 5596 34508
rect 5540 34372 5596 34428
rect 5540 34292 5596 34348
rect 8430 34532 8486 34588
rect 8430 34452 8486 34508
rect 8430 34372 8486 34428
rect 8430 34292 8486 34348
rect 11320 34532 11376 34588
rect 11320 34452 11376 34508
rect 11320 34372 11376 34428
rect 11320 34292 11376 34348
rect 14210 34532 14266 34588
rect 14210 34452 14266 34508
rect 14210 34372 14266 34428
rect 14210 34292 14266 34348
rect 17100 34532 17156 34588
rect 17100 34452 17156 34508
rect 17100 34372 17156 34428
rect 17100 34292 17156 34348
rect 19990 34532 20046 34588
rect 19990 34452 20046 34508
rect 19990 34372 20046 34428
rect 19990 34292 20046 34348
rect 22880 34532 22936 34588
rect 22880 34452 22936 34508
rect 22880 34372 22936 34428
rect 22880 34292 22936 34348
rect 25770 34532 25826 34588
rect 25770 34452 25826 34508
rect 25770 34372 25826 34428
rect 25770 34292 25826 34348
rect 28660 34532 28716 34588
rect 28660 34452 28716 34508
rect 28660 34372 28716 34428
rect 28660 34292 28716 34348
rect 31550 34532 31606 34588
rect 31550 34452 31606 34508
rect 31550 34372 31606 34428
rect 31550 34292 31606 34348
rect 34440 34532 34496 34588
rect 34440 34452 34496 34508
rect 34440 34372 34496 34428
rect 34440 34292 34496 34348
rect 37330 34532 37386 34588
rect 37330 34452 37386 34508
rect 37330 34372 37386 34428
rect 37330 34292 37386 34348
rect 40220 34532 40276 34588
rect 40220 34452 40276 34508
rect 40220 34372 40276 34428
rect 40220 34292 40276 34348
rect 43110 34532 43166 34588
rect 43110 34452 43166 34508
rect 43110 34372 43166 34428
rect 43110 34292 43166 34348
rect 46000 34532 46056 34588
rect 46000 34452 46056 34508
rect 46000 34372 46056 34428
rect 46000 34292 46056 34348
rect 49008 34532 49064 34588
rect 49008 34452 49064 34508
rect 49008 34372 49064 34428
rect 49008 34292 49064 34348
rect 52237 34532 52293 34588
rect 52237 34452 52293 34508
rect 52237 34372 52293 34428
rect 52237 34292 52293 34348
rect 53638 34532 53694 34588
rect 53638 34452 53694 34508
rect 53638 34372 53694 34428
rect 53638 34292 53694 34348
rect 53806 34532 53862 34588
rect 53806 34452 53862 34508
rect 53806 34372 53862 34428
rect 53806 34292 53862 34348
rect 54550 34532 54606 34588
rect 54550 34452 54606 34508
rect 54550 34372 54606 34428
rect 54550 34292 54606 34348
rect 54940 34532 54996 34588
rect 54940 34452 54996 34508
rect 54940 34372 54996 34428
rect 54940 34292 54996 34348
rect 55656 34532 55712 34588
rect 55656 34452 55712 34508
rect 55656 34372 55712 34428
rect 55656 34292 55712 34348
rect 56234 34532 56290 34588
rect 56234 34452 56290 34508
rect 56234 34372 56290 34428
rect 56234 34292 56290 34348
rect 56679 34532 56735 34588
rect 56679 34452 56735 34508
rect 56679 34372 56735 34428
rect 56679 34292 56735 34348
rect 56983 34532 57039 34588
rect 56983 34452 57039 34508
rect 56983 34372 57039 34428
rect 56983 34292 57039 34348
rect 57825 34532 57881 34588
rect 57825 34452 57881 34508
rect 57825 34372 57881 34428
rect 57825 34292 57881 34348
rect 58465 34532 58521 34588
rect 58465 34452 58521 34508
rect 58465 34372 58521 34428
rect 58465 34292 58521 34348
rect 59048 34532 59104 34588
rect 59048 34452 59104 34508
rect 59048 34372 59104 34428
rect 59048 34292 59104 34348
rect 60326 34532 60382 34588
rect 60326 34452 60382 34508
rect 60326 34372 60382 34428
rect 60326 34292 60382 34348
rect 60484 34532 60540 34588
rect 60484 34452 60540 34508
rect 60484 34372 60540 34428
rect 60484 34292 60540 34348
rect 62528 34532 62584 34588
rect 62608 34532 62664 34588
rect 62528 34452 62584 34508
rect 62608 34452 62664 34508
rect 62528 34372 62584 34428
rect 62608 34372 62664 34428
rect 62528 34292 62584 34348
rect 62608 34292 62664 34348
rect 2184 32180 2240 32236
rect 2264 32180 2320 32236
rect 2184 32100 2240 32156
rect 2264 32100 2320 32156
rect 2184 32020 2240 32076
rect 2264 32020 2320 32076
rect 2184 31940 2240 31996
rect 2264 31940 2320 31996
rect 5393 32180 5449 32236
rect 5393 32100 5449 32156
rect 5393 32020 5449 32076
rect 5393 31940 5449 31996
rect 8283 32180 8339 32236
rect 8283 32100 8339 32156
rect 8283 32020 8339 32076
rect 8283 31940 8339 31996
rect 11173 32180 11229 32236
rect 11173 32100 11229 32156
rect 11173 32020 11229 32076
rect 11173 31940 11229 31996
rect 14063 32180 14119 32236
rect 14063 32100 14119 32156
rect 14063 32020 14119 32076
rect 14063 31940 14119 31996
rect 16953 32180 17009 32236
rect 16953 32100 17009 32156
rect 16953 32020 17009 32076
rect 16953 31940 17009 31996
rect 19843 32180 19899 32236
rect 19843 32100 19899 32156
rect 19843 32020 19899 32076
rect 19843 31940 19899 31996
rect 22733 32180 22789 32236
rect 22733 32100 22789 32156
rect 22733 32020 22789 32076
rect 22733 31940 22789 31996
rect 25623 32180 25679 32236
rect 25623 32100 25679 32156
rect 25623 32020 25679 32076
rect 25623 31940 25679 31996
rect 28513 32180 28569 32236
rect 28513 32100 28569 32156
rect 28513 32020 28569 32076
rect 28513 31940 28569 31996
rect 31403 32180 31459 32236
rect 31403 32100 31459 32156
rect 31403 32020 31459 32076
rect 31403 31940 31459 31996
rect 34293 32180 34349 32236
rect 34293 32100 34349 32156
rect 34293 32020 34349 32076
rect 34293 31940 34349 31996
rect 37183 32180 37239 32236
rect 37183 32100 37239 32156
rect 37183 32020 37239 32076
rect 37183 31940 37239 31996
rect 40073 32180 40129 32236
rect 40073 32100 40129 32156
rect 40073 32020 40129 32076
rect 40073 31940 40129 31996
rect 42963 32180 43019 32236
rect 42963 32100 43019 32156
rect 42963 32020 43019 32076
rect 42963 31940 43019 31996
rect 45853 32180 45909 32236
rect 45853 32100 45909 32156
rect 45853 32020 45909 32076
rect 45853 31940 45909 31996
rect 48800 32180 48856 32236
rect 48800 32100 48856 32156
rect 48800 32020 48856 32076
rect 48800 31940 48856 31996
rect 49662 32180 49718 32236
rect 49742 32180 49798 32236
rect 49662 32100 49718 32156
rect 49742 32100 49798 32156
rect 49662 32020 49718 32076
rect 49742 32020 49798 32076
rect 49662 31940 49718 31996
rect 49742 31940 49798 31996
rect 52956 32180 53012 32236
rect 52956 32100 53012 32156
rect 52956 32020 53012 32076
rect 52956 31940 53012 31996
rect 53114 32180 53170 32236
rect 53114 32100 53170 32156
rect 53114 32020 53170 32076
rect 53114 31940 53170 31996
rect 53470 32180 53526 32236
rect 53470 32100 53526 32156
rect 53470 32020 53526 32076
rect 53470 31940 53526 31996
rect 54788 32180 54844 32236
rect 54788 32100 54844 32156
rect 54788 32020 54844 32076
rect 54788 31940 54844 31996
rect 55381 32180 55437 32236
rect 55381 32100 55437 32156
rect 55381 32020 55437 32076
rect 55381 31940 55437 31996
rect 56527 32180 56583 32236
rect 56527 32100 56583 32156
rect 56527 32020 56583 32076
rect 56527 31940 56583 31996
rect 57963 32180 58019 32236
rect 58043 32180 58099 32236
rect 57963 32100 58019 32156
rect 58043 32100 58099 32156
rect 57963 32020 58019 32076
rect 58043 32020 58099 32076
rect 57963 31940 58019 31996
rect 58043 31940 58099 31996
rect 59206 32180 59262 32236
rect 59206 32100 59262 32156
rect 59206 32020 59262 32076
rect 59206 31940 59262 31996
rect 59364 32180 59420 32236
rect 59364 32100 59420 32156
rect 59364 32020 59420 32076
rect 59364 31940 59420 31996
rect 59672 32180 59728 32236
rect 59672 32100 59728 32156
rect 59672 32020 59728 32076
rect 59672 31940 59728 31996
rect 59818 32180 59874 32236
rect 59818 32100 59874 32156
rect 59818 32020 59874 32076
rect 59818 31940 59874 31996
rect 59954 32180 60010 32236
rect 60034 32180 60090 32236
rect 59954 32100 60010 32156
rect 60034 32100 60090 32156
rect 59954 32020 60010 32076
rect 60034 32020 60090 32076
rect 59954 31940 60010 31996
rect 60034 31940 60090 31996
rect 62326 32180 62382 32236
rect 62406 32180 62462 32236
rect 62326 32100 62382 32156
rect 62406 32100 62462 32156
rect 62326 32020 62382 32076
rect 62406 32020 62462 32076
rect 62326 31940 62382 31996
rect 62406 31940 62462 31996
rect 2044 24532 2100 24588
rect 2044 24452 2100 24508
rect 2044 24372 2100 24428
rect 2044 24292 2100 24348
rect 5540 24532 5596 24588
rect 5540 24452 5596 24508
rect 5540 24372 5596 24428
rect 5540 24292 5596 24348
rect 8430 24532 8486 24588
rect 8430 24452 8486 24508
rect 8430 24372 8486 24428
rect 8430 24292 8486 24348
rect 11320 24532 11376 24588
rect 11320 24452 11376 24508
rect 11320 24372 11376 24428
rect 11320 24292 11376 24348
rect 14210 24532 14266 24588
rect 14210 24452 14266 24508
rect 14210 24372 14266 24428
rect 14210 24292 14266 24348
rect 17100 24532 17156 24588
rect 17100 24452 17156 24508
rect 17100 24372 17156 24428
rect 17100 24292 17156 24348
rect 19990 24532 20046 24588
rect 19990 24452 20046 24508
rect 19990 24372 20046 24428
rect 19990 24292 20046 24348
rect 22880 24532 22936 24588
rect 22880 24452 22936 24508
rect 22880 24372 22936 24428
rect 22880 24292 22936 24348
rect 25770 24532 25826 24588
rect 25770 24452 25826 24508
rect 25770 24372 25826 24428
rect 25770 24292 25826 24348
rect 28660 24532 28716 24588
rect 28660 24452 28716 24508
rect 28660 24372 28716 24428
rect 28660 24292 28716 24348
rect 31550 24532 31606 24588
rect 31550 24452 31606 24508
rect 31550 24372 31606 24428
rect 31550 24292 31606 24348
rect 34440 24532 34496 24588
rect 34440 24452 34496 24508
rect 34440 24372 34496 24428
rect 34440 24292 34496 24348
rect 37330 24532 37386 24588
rect 37330 24452 37386 24508
rect 37330 24372 37386 24428
rect 37330 24292 37386 24348
rect 40220 24532 40276 24588
rect 40220 24452 40276 24508
rect 40220 24372 40276 24428
rect 40220 24292 40276 24348
rect 43110 24532 43166 24588
rect 43110 24452 43166 24508
rect 43110 24372 43166 24428
rect 43110 24292 43166 24348
rect 46000 24532 46056 24588
rect 46000 24452 46056 24508
rect 46000 24372 46056 24428
rect 46000 24292 46056 24348
rect 49008 24532 49064 24588
rect 49008 24452 49064 24508
rect 49008 24372 49064 24428
rect 49008 24292 49064 24348
rect 52237 24532 52293 24588
rect 52237 24452 52293 24508
rect 52237 24372 52293 24428
rect 52237 24292 52293 24348
rect 53638 24532 53694 24588
rect 53638 24452 53694 24508
rect 53638 24372 53694 24428
rect 53638 24292 53694 24348
rect 53806 24532 53862 24588
rect 53806 24452 53862 24508
rect 53806 24372 53862 24428
rect 53806 24292 53862 24348
rect 54550 24532 54606 24588
rect 54550 24452 54606 24508
rect 54550 24372 54606 24428
rect 54550 24292 54606 24348
rect 54940 24532 54996 24588
rect 54940 24452 54996 24508
rect 54940 24372 54996 24428
rect 54940 24292 54996 24348
rect 55656 24532 55712 24588
rect 55656 24452 55712 24508
rect 55656 24372 55712 24428
rect 55656 24292 55712 24348
rect 56234 24532 56290 24588
rect 56234 24452 56290 24508
rect 56234 24372 56290 24428
rect 56234 24292 56290 24348
rect 56679 24532 56735 24588
rect 56679 24452 56735 24508
rect 56679 24372 56735 24428
rect 56679 24292 56735 24348
rect 56983 24532 57039 24588
rect 56983 24452 57039 24508
rect 56983 24372 57039 24428
rect 56983 24292 57039 24348
rect 57825 24532 57881 24588
rect 57825 24452 57881 24508
rect 57825 24372 57881 24428
rect 57825 24292 57881 24348
rect 58465 24532 58521 24588
rect 58465 24452 58521 24508
rect 58465 24372 58521 24428
rect 58465 24292 58521 24348
rect 59048 24532 59104 24588
rect 59048 24452 59104 24508
rect 59048 24372 59104 24428
rect 59048 24292 59104 24348
rect 60326 24532 60382 24588
rect 60326 24452 60382 24508
rect 60326 24372 60382 24428
rect 60326 24292 60382 24348
rect 60484 24532 60540 24588
rect 60484 24452 60540 24508
rect 60484 24372 60540 24428
rect 60484 24292 60540 24348
rect 62528 24532 62584 24588
rect 62608 24532 62664 24588
rect 62528 24452 62584 24508
rect 62608 24452 62664 24508
rect 62528 24372 62584 24428
rect 62608 24372 62664 24428
rect 62528 24292 62584 24348
rect 62608 24292 62664 24348
rect 2184 22180 2240 22236
rect 2264 22180 2320 22236
rect 2184 22100 2240 22156
rect 2264 22100 2320 22156
rect 2184 22020 2240 22076
rect 2264 22020 2320 22076
rect 2184 21940 2240 21996
rect 2264 21940 2320 21996
rect 5393 22180 5449 22236
rect 5393 22100 5449 22156
rect 5393 22020 5449 22076
rect 5393 21940 5449 21996
rect 8283 22180 8339 22236
rect 8283 22100 8339 22156
rect 8283 22020 8339 22076
rect 8283 21940 8339 21996
rect 11173 22180 11229 22236
rect 11173 22100 11229 22156
rect 11173 22020 11229 22076
rect 11173 21940 11229 21996
rect 14063 22180 14119 22236
rect 14063 22100 14119 22156
rect 14063 22020 14119 22076
rect 14063 21940 14119 21996
rect 16953 22180 17009 22236
rect 16953 22100 17009 22156
rect 16953 22020 17009 22076
rect 16953 21940 17009 21996
rect 19843 22180 19899 22236
rect 19843 22100 19899 22156
rect 19843 22020 19899 22076
rect 19843 21940 19899 21996
rect 22733 22180 22789 22236
rect 22733 22100 22789 22156
rect 22733 22020 22789 22076
rect 22733 21940 22789 21996
rect 25623 22180 25679 22236
rect 25623 22100 25679 22156
rect 25623 22020 25679 22076
rect 25623 21940 25679 21996
rect 28513 22180 28569 22236
rect 28513 22100 28569 22156
rect 28513 22020 28569 22076
rect 28513 21940 28569 21996
rect 31403 22180 31459 22236
rect 31403 22100 31459 22156
rect 31403 22020 31459 22076
rect 31403 21940 31459 21996
rect 34293 22180 34349 22236
rect 34293 22100 34349 22156
rect 34293 22020 34349 22076
rect 34293 21940 34349 21996
rect 37183 22180 37239 22236
rect 37183 22100 37239 22156
rect 37183 22020 37239 22076
rect 37183 21940 37239 21996
rect 40073 22180 40129 22236
rect 40073 22100 40129 22156
rect 40073 22020 40129 22076
rect 40073 21940 40129 21996
rect 42963 22180 43019 22236
rect 42963 22100 43019 22156
rect 42963 22020 43019 22076
rect 42963 21940 43019 21996
rect 45853 22180 45909 22236
rect 45853 22100 45909 22156
rect 45853 22020 45909 22076
rect 45853 21940 45909 21996
rect 48800 22180 48856 22236
rect 48800 22100 48856 22156
rect 48800 22020 48856 22076
rect 48800 21940 48856 21996
rect 49662 22180 49718 22236
rect 49742 22180 49798 22236
rect 49662 22100 49718 22156
rect 49742 22100 49798 22156
rect 49662 22020 49718 22076
rect 49742 22020 49798 22076
rect 49662 21940 49718 21996
rect 49742 21940 49798 21996
rect 52956 22180 53012 22236
rect 52956 22100 53012 22156
rect 52956 22020 53012 22076
rect 52956 21940 53012 21996
rect 53114 22180 53170 22236
rect 53114 22100 53170 22156
rect 53114 22020 53170 22076
rect 53114 21940 53170 21996
rect 53470 22180 53526 22236
rect 53470 22100 53526 22156
rect 53470 22020 53526 22076
rect 53470 21940 53526 21996
rect 54788 22180 54844 22236
rect 54788 22100 54844 22156
rect 54788 22020 54844 22076
rect 54788 21940 54844 21996
rect 55381 22180 55437 22236
rect 55381 22100 55437 22156
rect 55381 22020 55437 22076
rect 55381 21940 55437 21996
rect 56527 22180 56583 22236
rect 56527 22100 56583 22156
rect 56527 22020 56583 22076
rect 56527 21940 56583 21996
rect 57963 22180 58019 22236
rect 58043 22180 58099 22236
rect 57963 22100 58019 22156
rect 58043 22100 58099 22156
rect 57963 22020 58019 22076
rect 58043 22020 58099 22076
rect 57963 21940 58019 21996
rect 58043 21940 58099 21996
rect 59206 22180 59262 22236
rect 59206 22100 59262 22156
rect 59206 22020 59262 22076
rect 59206 21940 59262 21996
rect 59364 22180 59420 22236
rect 59364 22100 59420 22156
rect 59364 22020 59420 22076
rect 59364 21940 59420 21996
rect 59672 22180 59728 22236
rect 59672 22100 59728 22156
rect 59672 22020 59728 22076
rect 59672 21940 59728 21996
rect 59818 22180 59874 22236
rect 59818 22100 59874 22156
rect 59818 22020 59874 22076
rect 59818 21940 59874 21996
rect 59954 22180 60010 22236
rect 60034 22180 60090 22236
rect 59954 22100 60010 22156
rect 60034 22100 60090 22156
rect 59954 22020 60010 22076
rect 60034 22020 60090 22076
rect 59954 21940 60010 21996
rect 60034 21940 60090 21996
rect 62326 22180 62382 22236
rect 62406 22180 62462 22236
rect 62326 22100 62382 22156
rect 62406 22100 62462 22156
rect 62326 22020 62382 22076
rect 62406 22020 62462 22076
rect 62326 21940 62382 21996
rect 62406 21940 62462 21996
rect 2044 14532 2100 14588
rect 2044 14452 2100 14508
rect 2044 14372 2100 14428
rect 2044 14292 2100 14348
rect 5540 14532 5596 14588
rect 5540 14452 5596 14508
rect 5540 14372 5596 14428
rect 5540 14292 5596 14348
rect 8430 14532 8486 14588
rect 8430 14452 8486 14508
rect 8430 14372 8486 14428
rect 8430 14292 8486 14348
rect 11320 14532 11376 14588
rect 11320 14452 11376 14508
rect 11320 14372 11376 14428
rect 11320 14292 11376 14348
rect 14210 14532 14266 14588
rect 14210 14452 14266 14508
rect 14210 14372 14266 14428
rect 14210 14292 14266 14348
rect 17100 14532 17156 14588
rect 17100 14452 17156 14508
rect 17100 14372 17156 14428
rect 17100 14292 17156 14348
rect 19990 14532 20046 14588
rect 19990 14452 20046 14508
rect 19990 14372 20046 14428
rect 19990 14292 20046 14348
rect 22880 14532 22936 14588
rect 22880 14452 22936 14508
rect 22880 14372 22936 14428
rect 22880 14292 22936 14348
rect 25770 14532 25826 14588
rect 25770 14452 25826 14508
rect 25770 14372 25826 14428
rect 25770 14292 25826 14348
rect 28660 14532 28716 14588
rect 28660 14452 28716 14508
rect 28660 14372 28716 14428
rect 28660 14292 28716 14348
rect 31550 14532 31606 14588
rect 31550 14452 31606 14508
rect 31550 14372 31606 14428
rect 31550 14292 31606 14348
rect 34440 14532 34496 14588
rect 34440 14452 34496 14508
rect 34440 14372 34496 14428
rect 34440 14292 34496 14348
rect 37330 14532 37386 14588
rect 37330 14452 37386 14508
rect 37330 14372 37386 14428
rect 37330 14292 37386 14348
rect 40220 14532 40276 14588
rect 40220 14452 40276 14508
rect 40220 14372 40276 14428
rect 40220 14292 40276 14348
rect 43110 14532 43166 14588
rect 43110 14452 43166 14508
rect 43110 14372 43166 14428
rect 43110 14292 43166 14348
rect 46000 14532 46056 14588
rect 46000 14452 46056 14508
rect 46000 14372 46056 14428
rect 46000 14292 46056 14348
rect 49008 14532 49064 14588
rect 49008 14452 49064 14508
rect 49008 14372 49064 14428
rect 49008 14292 49064 14348
rect 52237 14532 52293 14588
rect 52237 14452 52293 14508
rect 52237 14372 52293 14428
rect 52237 14292 52293 14348
rect 53638 14532 53694 14588
rect 53638 14452 53694 14508
rect 53638 14372 53694 14428
rect 53638 14292 53694 14348
rect 53806 14532 53862 14588
rect 53806 14452 53862 14508
rect 53806 14372 53862 14428
rect 53806 14292 53862 14348
rect 54550 14532 54606 14588
rect 54550 14452 54606 14508
rect 54550 14372 54606 14428
rect 54550 14292 54606 14348
rect 54940 14532 54996 14588
rect 54940 14452 54996 14508
rect 54940 14372 54996 14428
rect 54940 14292 54996 14348
rect 55656 14532 55712 14588
rect 55656 14452 55712 14508
rect 55656 14372 55712 14428
rect 55656 14292 55712 14348
rect 56234 14532 56290 14588
rect 56234 14452 56290 14508
rect 56234 14372 56290 14428
rect 56234 14292 56290 14348
rect 56679 14532 56735 14588
rect 56679 14452 56735 14508
rect 56679 14372 56735 14428
rect 56679 14292 56735 14348
rect 56983 14532 57039 14588
rect 56983 14452 57039 14508
rect 56983 14372 57039 14428
rect 56983 14292 57039 14348
rect 57825 14532 57881 14588
rect 57825 14452 57881 14508
rect 57825 14372 57881 14428
rect 57825 14292 57881 14348
rect 58465 14532 58521 14588
rect 58465 14452 58521 14508
rect 58465 14372 58521 14428
rect 58465 14292 58521 14348
rect 59048 14532 59104 14588
rect 59048 14452 59104 14508
rect 59048 14372 59104 14428
rect 59048 14292 59104 14348
rect 60326 14532 60382 14588
rect 60326 14452 60382 14508
rect 60326 14372 60382 14428
rect 60326 14292 60382 14348
rect 60484 14532 60540 14588
rect 60484 14452 60540 14508
rect 60484 14372 60540 14428
rect 60484 14292 60540 14348
rect 62528 14532 62584 14588
rect 62608 14532 62664 14588
rect 62528 14452 62584 14508
rect 62608 14452 62664 14508
rect 62528 14372 62584 14428
rect 62608 14372 62664 14428
rect 62528 14292 62584 14348
rect 62608 14292 62664 14348
rect 2184 12180 2240 12236
rect 2264 12180 2320 12236
rect 2184 12100 2240 12156
rect 2264 12100 2320 12156
rect 2184 12020 2240 12076
rect 2264 12020 2320 12076
rect 2184 11940 2240 11996
rect 2264 11940 2320 11996
rect 5393 12180 5449 12236
rect 5393 12100 5449 12156
rect 5393 12020 5449 12076
rect 5393 11940 5449 11996
rect 8283 12180 8339 12236
rect 8283 12100 8339 12156
rect 8283 12020 8339 12076
rect 8283 11940 8339 11996
rect 11173 12180 11229 12236
rect 11173 12100 11229 12156
rect 11173 12020 11229 12076
rect 11173 11940 11229 11996
rect 14063 12180 14119 12236
rect 14063 12100 14119 12156
rect 14063 12020 14119 12076
rect 14063 11940 14119 11996
rect 16953 12180 17009 12236
rect 16953 12100 17009 12156
rect 16953 12020 17009 12076
rect 16953 11940 17009 11996
rect 19843 12180 19899 12236
rect 19843 12100 19899 12156
rect 19843 12020 19899 12076
rect 19843 11940 19899 11996
rect 22733 12180 22789 12236
rect 22733 12100 22789 12156
rect 22733 12020 22789 12076
rect 22733 11940 22789 11996
rect 25623 12180 25679 12236
rect 25623 12100 25679 12156
rect 25623 12020 25679 12076
rect 25623 11940 25679 11996
rect 28513 12180 28569 12236
rect 28513 12100 28569 12156
rect 28513 12020 28569 12076
rect 28513 11940 28569 11996
rect 31403 12180 31459 12236
rect 31403 12100 31459 12156
rect 31403 12020 31459 12076
rect 31403 11940 31459 11996
rect 34293 12180 34349 12236
rect 34293 12100 34349 12156
rect 34293 12020 34349 12076
rect 34293 11940 34349 11996
rect 37183 12180 37239 12236
rect 37183 12100 37239 12156
rect 37183 12020 37239 12076
rect 37183 11940 37239 11996
rect 40073 12180 40129 12236
rect 40073 12100 40129 12156
rect 40073 12020 40129 12076
rect 40073 11940 40129 11996
rect 42963 12180 43019 12236
rect 42963 12100 43019 12156
rect 42963 12020 43019 12076
rect 42963 11940 43019 11996
rect 45853 12180 45909 12236
rect 45853 12100 45909 12156
rect 45853 12020 45909 12076
rect 45853 11940 45909 11996
rect 48800 12180 48856 12236
rect 48800 12100 48856 12156
rect 48800 12020 48856 12076
rect 48800 11940 48856 11996
rect 49662 12180 49718 12236
rect 49742 12180 49798 12236
rect 49662 12100 49718 12156
rect 49742 12100 49798 12156
rect 49662 12020 49718 12076
rect 49742 12020 49798 12076
rect 49662 11940 49718 11996
rect 49742 11940 49798 11996
rect 52956 12180 53012 12236
rect 52956 12100 53012 12156
rect 52956 12020 53012 12076
rect 52956 11940 53012 11996
rect 53114 12180 53170 12236
rect 53114 12100 53170 12156
rect 53114 12020 53170 12076
rect 53114 11940 53170 11996
rect 53470 12180 53526 12236
rect 53470 12100 53526 12156
rect 53470 12020 53526 12076
rect 53470 11940 53526 11996
rect 54788 12180 54844 12236
rect 54788 12100 54844 12156
rect 54788 12020 54844 12076
rect 54788 11940 54844 11996
rect 55381 12180 55437 12236
rect 55381 12100 55437 12156
rect 55381 12020 55437 12076
rect 55381 11940 55437 11996
rect 56527 12180 56583 12236
rect 56527 12100 56583 12156
rect 56527 12020 56583 12076
rect 56527 11940 56583 11996
rect 57963 12180 58019 12236
rect 58043 12180 58099 12236
rect 57963 12100 58019 12156
rect 58043 12100 58099 12156
rect 57963 12020 58019 12076
rect 58043 12020 58099 12076
rect 57963 11940 58019 11996
rect 58043 11940 58099 11996
rect 59206 12180 59262 12236
rect 59206 12100 59262 12156
rect 59206 12020 59262 12076
rect 59206 11940 59262 11996
rect 59364 12180 59420 12236
rect 59364 12100 59420 12156
rect 59364 12020 59420 12076
rect 59364 11940 59420 11996
rect 59672 12180 59728 12236
rect 59672 12100 59728 12156
rect 59672 12020 59728 12076
rect 59672 11940 59728 11996
rect 59818 12180 59874 12236
rect 59818 12100 59874 12156
rect 59818 12020 59874 12076
rect 59818 11940 59874 11996
rect 59954 12180 60010 12236
rect 60034 12180 60090 12236
rect 59954 12100 60010 12156
rect 60034 12100 60090 12156
rect 59954 12020 60010 12076
rect 60034 12020 60090 12076
rect 59954 11940 60010 11996
rect 60034 11940 60090 11996
rect 62326 12180 62382 12236
rect 62406 12180 62462 12236
rect 62326 12100 62382 12156
rect 62406 12100 62462 12156
rect 62326 12020 62382 12076
rect 62406 12020 62462 12076
rect 62326 11940 62382 11996
rect 62406 11940 62462 11996
rect 30838 7656 30894 7712
rect 30286 7520 30342 7576
rect 1864 2180 1920 2236
rect 1944 2180 2000 2236
rect 2024 2180 2080 2236
rect 2104 2180 2160 2236
rect 1864 2100 1920 2156
rect 1944 2100 2000 2156
rect 2024 2100 2080 2156
rect 2104 2100 2160 2156
rect 1864 2020 1920 2076
rect 1944 2020 2000 2076
rect 2024 2020 2080 2076
rect 2104 2020 2160 2076
rect 1864 1940 1920 1996
rect 1944 1940 2000 1996
rect 2024 1940 2080 1996
rect 2104 1940 2160 1996
rect 4216 4532 4272 4588
rect 4296 4532 4352 4588
rect 4376 4532 4432 4588
rect 4456 4532 4512 4588
rect 4216 4452 4272 4508
rect 4296 4452 4352 4508
rect 4376 4452 4432 4508
rect 4456 4452 4512 4508
rect 4216 4378 4272 4428
rect 4296 4378 4352 4428
rect 4376 4378 4432 4428
rect 4456 4378 4512 4428
rect 4216 4372 4262 4378
rect 4262 4372 4272 4378
rect 4296 4372 4326 4378
rect 4326 4372 4338 4378
rect 4338 4372 4352 4378
rect 4376 4372 4390 4378
rect 4390 4372 4402 4378
rect 4402 4372 4432 4378
rect 4456 4372 4466 4378
rect 4466 4372 4512 4378
rect 4216 4326 4262 4348
rect 4262 4326 4272 4348
rect 4296 4326 4326 4348
rect 4326 4326 4338 4348
rect 4338 4326 4352 4348
rect 4376 4326 4390 4348
rect 4390 4326 4402 4348
rect 4402 4326 4432 4348
rect 4456 4326 4466 4348
rect 4466 4326 4512 4348
rect 4216 4292 4272 4326
rect 4296 4292 4352 4326
rect 4376 4292 4432 4326
rect 4456 4292 4512 4326
rect 11864 2180 11920 2236
rect 11944 2180 12000 2236
rect 12024 2180 12080 2236
rect 12104 2180 12160 2236
rect 11864 2100 11920 2156
rect 11944 2100 12000 2156
rect 12024 2100 12080 2156
rect 12104 2100 12160 2156
rect 11864 2020 11920 2076
rect 11944 2020 12000 2076
rect 12024 2020 12080 2076
rect 12104 2020 12160 2076
rect 11864 1940 11920 1996
rect 11944 1940 12000 1996
rect 12024 1940 12080 1996
rect 12104 1940 12160 1996
rect 14216 4532 14272 4588
rect 14296 4532 14352 4588
rect 14376 4532 14432 4588
rect 14456 4532 14512 4588
rect 14216 4452 14272 4508
rect 14296 4452 14352 4508
rect 14376 4452 14432 4508
rect 14456 4452 14512 4508
rect 14216 4378 14272 4428
rect 14296 4378 14352 4428
rect 14376 4378 14432 4428
rect 14456 4378 14512 4428
rect 14216 4372 14262 4378
rect 14262 4372 14272 4378
rect 14296 4372 14326 4378
rect 14326 4372 14338 4378
rect 14338 4372 14352 4378
rect 14376 4372 14390 4378
rect 14390 4372 14402 4378
rect 14402 4372 14432 4378
rect 14456 4372 14466 4378
rect 14466 4372 14512 4378
rect 14216 4326 14262 4348
rect 14262 4326 14272 4348
rect 14296 4326 14326 4348
rect 14326 4326 14338 4348
rect 14338 4326 14352 4348
rect 14376 4326 14390 4348
rect 14390 4326 14402 4348
rect 14402 4326 14432 4348
rect 14456 4326 14466 4348
rect 14466 4326 14512 4348
rect 14216 4292 14272 4326
rect 14296 4292 14352 4326
rect 14376 4292 14432 4326
rect 14456 4292 14512 4326
rect 24582 5888 24638 5944
rect 14738 3304 14794 3360
rect 20902 3188 20958 3224
rect 20902 3168 20904 3188
rect 20904 3168 20956 3188
rect 20956 3168 20958 3188
rect 21864 2180 21920 2236
rect 21944 2180 22000 2236
rect 22024 2180 22080 2236
rect 22104 2180 22160 2236
rect 21864 2100 21920 2156
rect 21944 2100 22000 2156
rect 22024 2100 22080 2156
rect 22104 2100 22160 2156
rect 21864 2020 21920 2076
rect 21944 2020 22000 2076
rect 22024 2020 22080 2076
rect 22104 2020 22160 2076
rect 21864 1940 21920 1996
rect 21944 1940 22000 1996
rect 22024 1940 22080 1996
rect 22104 1940 22160 1996
rect 23202 1400 23258 1456
rect 24216 4532 24272 4588
rect 24296 4532 24352 4588
rect 24376 4532 24432 4588
rect 24456 4532 24512 4588
rect 24216 4452 24272 4508
rect 24296 4452 24352 4508
rect 24376 4452 24432 4508
rect 24456 4452 24512 4508
rect 24216 4378 24272 4428
rect 24296 4378 24352 4428
rect 24376 4378 24432 4428
rect 24456 4378 24512 4428
rect 24216 4372 24262 4378
rect 24262 4372 24272 4378
rect 24296 4372 24326 4378
rect 24326 4372 24338 4378
rect 24338 4372 24352 4378
rect 24376 4372 24390 4378
rect 24390 4372 24402 4378
rect 24402 4372 24432 4378
rect 24456 4372 24466 4378
rect 24466 4372 24512 4378
rect 24216 4326 24262 4348
rect 24262 4326 24272 4348
rect 24296 4326 24326 4348
rect 24326 4326 24338 4348
rect 24338 4326 24352 4348
rect 24376 4326 24390 4348
rect 24390 4326 24402 4348
rect 24402 4326 24432 4348
rect 24456 4326 24466 4348
rect 24466 4326 24512 4348
rect 24216 4292 24272 4326
rect 24296 4292 24352 4326
rect 24376 4292 24432 4326
rect 24456 4292 24512 4326
rect 25778 5092 25834 5128
rect 25778 5072 25780 5092
rect 25780 5072 25832 5092
rect 25832 5072 25834 5092
rect 25870 3168 25926 3224
rect 26146 3032 26202 3088
rect 27158 5208 27214 5264
rect 29090 6704 29146 6760
rect 28446 6432 28502 6488
rect 28078 5072 28134 5128
rect 27802 4936 27858 4992
rect 29734 6568 29790 6624
rect 28906 3052 28962 3088
rect 28906 3032 28908 3052
rect 28908 3032 28960 3052
rect 28960 3032 28962 3052
rect 41050 6840 41106 6896
rect 29734 4936 29790 4992
rect 28446 1420 28502 1456
rect 28446 1400 28448 1420
rect 28448 1400 28500 1420
rect 28500 1400 28502 1420
rect 31298 3984 31354 4040
rect 31114 1536 31170 1592
rect 32218 3032 32274 3088
rect 31864 2180 31920 2236
rect 31944 2180 32000 2236
rect 32024 2180 32080 2236
rect 32104 2180 32160 2236
rect 31864 2100 31920 2156
rect 31944 2100 32000 2156
rect 32024 2100 32080 2156
rect 32104 2100 32160 2156
rect 31864 2020 31920 2076
rect 31944 2020 32000 2076
rect 32024 2020 32080 2076
rect 32104 2020 32160 2076
rect 31864 1940 31920 1996
rect 31944 1940 32000 1996
rect 32024 1940 32080 1996
rect 32104 1940 32160 1996
rect 34058 4800 34114 4856
rect 34216 4532 34272 4588
rect 34296 4532 34352 4588
rect 34376 4532 34432 4588
rect 34456 4532 34512 4588
rect 34216 4452 34272 4508
rect 34296 4452 34352 4508
rect 34376 4452 34432 4508
rect 34456 4452 34512 4508
rect 34216 4378 34272 4428
rect 34296 4378 34352 4428
rect 34376 4378 34432 4428
rect 34456 4378 34512 4428
rect 34216 4372 34262 4378
rect 34262 4372 34272 4378
rect 34296 4372 34326 4378
rect 34326 4372 34338 4378
rect 34338 4372 34352 4378
rect 34376 4372 34390 4378
rect 34390 4372 34402 4378
rect 34402 4372 34432 4378
rect 34456 4372 34466 4378
rect 34466 4372 34512 4378
rect 34216 4326 34262 4348
rect 34262 4326 34272 4348
rect 34296 4326 34326 4348
rect 34326 4326 34338 4348
rect 34338 4326 34352 4348
rect 34376 4326 34390 4348
rect 34390 4326 34402 4348
rect 34402 4326 34432 4348
rect 34456 4326 34466 4348
rect 34466 4326 34512 4348
rect 34216 4292 34272 4326
rect 34296 4292 34352 4326
rect 34376 4292 34432 4326
rect 34456 4292 34512 4326
rect 40406 5752 40462 5808
rect 37002 5636 37058 5672
rect 37002 5616 37004 5636
rect 37004 5616 37056 5636
rect 37056 5616 37058 5636
rect 44638 6024 44694 6080
rect 35990 1536 36046 1592
rect 41418 3304 41474 3360
rect 41694 5616 41750 5672
rect 42706 5108 42708 5128
rect 42708 5108 42760 5128
rect 42760 5108 42762 5128
rect 42706 5072 42762 5108
rect 43350 4120 43406 4176
rect 41864 2180 41920 2236
rect 41944 2180 42000 2236
rect 42024 2180 42080 2236
rect 42104 2180 42160 2236
rect 41864 2100 41920 2156
rect 41944 2100 42000 2156
rect 42024 2100 42080 2156
rect 42104 2100 42160 2156
rect 41864 2020 41920 2076
rect 41944 2020 42000 2076
rect 42024 2020 42080 2076
rect 42104 2020 42160 2076
rect 41864 1940 41920 1996
rect 41944 1940 42000 1996
rect 42024 1940 42080 1996
rect 42104 1940 42160 1996
rect 46754 6160 46810 6216
rect 46202 5344 46258 5400
rect 44216 4532 44272 4588
rect 44296 4532 44352 4588
rect 44376 4532 44432 4588
rect 44456 4532 44512 4588
rect 44216 4452 44272 4508
rect 44296 4452 44352 4508
rect 44376 4452 44432 4508
rect 44456 4452 44512 4508
rect 44216 4378 44272 4428
rect 44296 4378 44352 4428
rect 44376 4378 44432 4428
rect 44456 4378 44512 4428
rect 44216 4372 44262 4378
rect 44262 4372 44272 4378
rect 44296 4372 44326 4378
rect 44326 4372 44338 4378
rect 44338 4372 44352 4378
rect 44376 4372 44390 4378
rect 44390 4372 44402 4378
rect 44402 4372 44432 4378
rect 44456 4372 44466 4378
rect 44466 4372 44512 4378
rect 44216 4326 44262 4348
rect 44262 4326 44272 4348
rect 44296 4326 44326 4348
rect 44326 4326 44338 4348
rect 44338 4326 44352 4348
rect 44376 4326 44390 4348
rect 44390 4326 44402 4348
rect 44402 4326 44432 4348
rect 44456 4326 44466 4348
rect 44466 4326 44512 4348
rect 44216 4292 44272 4326
rect 44296 4292 44352 4326
rect 44376 4292 44432 4326
rect 44456 4292 44512 4326
rect 44730 4936 44786 4992
rect 44730 4120 44786 4176
rect 48962 5480 49018 5536
rect 51864 2180 51920 2236
rect 51944 2180 52000 2236
rect 52024 2180 52080 2236
rect 52104 2180 52160 2236
rect 51864 2100 51920 2156
rect 51944 2100 52000 2156
rect 52024 2100 52080 2156
rect 52104 2100 52160 2156
rect 51864 2020 51920 2076
rect 51944 2020 52000 2076
rect 52024 2020 52080 2076
rect 52104 2020 52160 2076
rect 51864 1940 51920 1996
rect 51944 1940 52000 1996
rect 52024 1940 52080 1996
rect 52104 1940 52160 1996
rect 55862 6296 55918 6352
rect 55862 6024 55918 6080
rect 54216 4532 54272 4588
rect 54296 4532 54352 4588
rect 54376 4532 54432 4588
rect 54456 4532 54512 4588
rect 54216 4452 54272 4508
rect 54296 4452 54352 4508
rect 54376 4452 54432 4508
rect 54456 4452 54512 4508
rect 54216 4378 54272 4428
rect 54296 4378 54352 4428
rect 54376 4378 54432 4428
rect 54456 4378 54512 4428
rect 54216 4372 54262 4378
rect 54262 4372 54272 4378
rect 54296 4372 54326 4378
rect 54326 4372 54338 4378
rect 54338 4372 54352 4378
rect 54376 4372 54390 4378
rect 54390 4372 54402 4378
rect 54402 4372 54432 4378
rect 54456 4372 54466 4378
rect 54466 4372 54512 4378
rect 54216 4326 54262 4348
rect 54262 4326 54272 4348
rect 54296 4326 54326 4348
rect 54326 4326 54338 4348
rect 54338 4326 54352 4348
rect 54376 4326 54390 4348
rect 54390 4326 54402 4348
rect 54402 4326 54432 4348
rect 54456 4326 54466 4348
rect 54466 4326 54512 4348
rect 54216 4292 54272 4326
rect 54296 4292 54352 4326
rect 54376 4292 54432 4326
rect 54456 4292 54512 4326
rect 55954 5480 56010 5536
rect 58162 5888 58218 5944
rect 59726 6024 59782 6080
rect 61566 6976 61622 7032
rect 61014 5480 61070 5536
rect 61566 5752 61622 5808
rect 62302 6568 62358 6624
rect 63774 52536 63830 52592
rect 63774 50260 63776 50280
rect 63776 50260 63828 50280
rect 63828 50260 63830 50280
rect 63774 50224 63830 50260
rect 64970 48084 64972 48104
rect 64972 48084 65024 48104
rect 65024 48084 65026 48104
rect 64970 48048 65026 48084
rect 64418 47676 64420 47696
rect 64420 47676 64472 47696
rect 64472 47676 64474 47696
rect 64418 47640 64474 47676
rect 63774 43308 63830 43344
rect 63774 43288 63776 43308
rect 63776 43288 63828 43308
rect 63828 43288 63830 43308
rect 63682 17856 63738 17912
rect 63682 11736 63738 11792
rect 61750 6160 61806 6216
rect 62302 6160 62358 6216
rect 61750 5752 61806 5808
rect 60646 4120 60702 4176
rect 62946 6840 63002 6896
rect 62762 5888 62818 5944
rect 61382 4120 61438 4176
rect 63406 5516 63408 5536
rect 63408 5516 63460 5536
rect 63460 5516 63462 5536
rect 63406 5480 63462 5516
rect 63314 5208 63370 5264
rect 63958 6296 64014 6352
rect 64694 12416 64750 12472
rect 63590 5208 63646 5264
rect 64970 7656 65026 7712
rect 64216 4532 64272 4588
rect 64296 4532 64352 4588
rect 64376 4532 64432 4588
rect 64456 4532 64512 4588
rect 64216 4452 64272 4508
rect 64296 4452 64352 4508
rect 64376 4452 64432 4508
rect 64456 4452 64512 4508
rect 64216 4378 64272 4428
rect 64296 4378 64352 4428
rect 64376 4378 64432 4428
rect 64456 4378 64512 4428
rect 64216 4372 64262 4378
rect 64262 4372 64272 4378
rect 64296 4372 64326 4378
rect 64326 4372 64338 4378
rect 64338 4372 64352 4378
rect 64376 4372 64390 4378
rect 64390 4372 64402 4378
rect 64402 4372 64432 4378
rect 64456 4372 64466 4378
rect 64466 4372 64512 4378
rect 64216 4326 64262 4348
rect 64262 4326 64272 4348
rect 64296 4326 64326 4348
rect 64326 4326 64338 4348
rect 64338 4326 64352 4348
rect 64376 4326 64390 4348
rect 64390 4326 64402 4348
rect 64402 4326 64432 4348
rect 64456 4326 64466 4348
rect 64466 4326 64512 4348
rect 64216 4292 64272 4326
rect 64296 4292 64352 4326
rect 64376 4292 64432 4326
rect 64456 4292 64512 4326
rect 63590 3032 63646 3088
rect 61864 2180 61920 2236
rect 61944 2180 62000 2236
rect 62024 2180 62080 2236
rect 62104 2180 62160 2236
rect 61864 2100 61920 2156
rect 61944 2100 62000 2156
rect 62024 2100 62080 2156
rect 62104 2100 62160 2156
rect 61864 2020 61920 2076
rect 61944 2020 62000 2076
rect 62024 2020 62080 2076
rect 62104 2020 62160 2076
rect 61864 1940 61920 1996
rect 61944 1940 62000 1996
rect 62024 1940 62080 1996
rect 62104 1940 62160 1996
rect 64878 5072 64934 5128
rect 65246 44784 65302 44840
rect 65246 40840 65302 40896
rect 65246 38664 65302 38720
rect 65614 33224 65670 33280
rect 65522 19116 65524 19136
rect 65524 19116 65576 19136
rect 65576 19116 65578 19136
rect 65522 19080 65578 19116
rect 65430 11464 65486 11520
rect 65246 6432 65302 6488
rect 65706 6568 65762 6624
rect 65982 5752 66038 5808
rect 66350 23432 66406 23488
rect 66350 23296 66406 23352
rect 66534 23432 66590 23488
rect 66994 23840 67050 23896
rect 71864 82180 71920 82236
rect 71944 82180 72000 82236
rect 72024 82180 72080 82236
rect 72104 82180 72160 82236
rect 71864 82118 71910 82156
rect 71910 82118 71920 82156
rect 71944 82118 71974 82156
rect 71974 82118 71986 82156
rect 71986 82118 72000 82156
rect 72024 82118 72038 82156
rect 72038 82118 72050 82156
rect 72050 82118 72080 82156
rect 72104 82118 72114 82156
rect 72114 82118 72160 82156
rect 71864 82100 71920 82118
rect 71944 82100 72000 82118
rect 72024 82100 72080 82118
rect 72104 82100 72160 82118
rect 71864 82020 71920 82076
rect 71944 82020 72000 82076
rect 72024 82020 72080 82076
rect 72104 82020 72160 82076
rect 71864 81940 71920 81996
rect 71944 81940 72000 81996
rect 72024 81940 72080 81996
rect 72104 81940 72160 81996
rect 71864 72180 71920 72236
rect 71944 72180 72000 72236
rect 72024 72180 72080 72236
rect 72104 72180 72160 72236
rect 71864 72100 71920 72156
rect 71944 72100 72000 72156
rect 72024 72100 72080 72156
rect 72104 72100 72160 72156
rect 71864 72020 71920 72076
rect 71944 72020 72000 72076
rect 72024 72020 72080 72076
rect 72104 72020 72160 72076
rect 71864 71940 71920 71996
rect 71944 71940 72000 71996
rect 72024 71940 72080 71996
rect 72104 71940 72160 71996
rect 71864 62180 71920 62236
rect 71944 62180 72000 62236
rect 72024 62180 72080 62236
rect 72104 62180 72160 62236
rect 71864 62100 71920 62156
rect 71944 62100 72000 62156
rect 72024 62100 72080 62156
rect 72104 62100 72160 62156
rect 71864 62020 71920 62076
rect 71944 62020 72000 62076
rect 72024 62020 72080 62076
rect 72104 62020 72160 62076
rect 71864 61940 71920 61996
rect 71944 61940 72000 61996
rect 72024 61940 72080 61996
rect 72104 61940 72160 61996
rect 70398 6024 70454 6080
rect 71864 52180 71920 52236
rect 71944 52180 72000 52236
rect 72024 52180 72080 52236
rect 72104 52180 72160 52236
rect 71864 52100 71920 52156
rect 71944 52100 72000 52156
rect 72024 52100 72080 52156
rect 72104 52100 72160 52156
rect 71864 52020 71920 52076
rect 71944 52020 72000 52076
rect 72024 52020 72080 52076
rect 72104 52020 72160 52076
rect 71864 51940 71920 51996
rect 71944 51940 72000 51996
rect 72024 51940 72080 51996
rect 72104 51940 72160 51996
rect 71864 42180 71920 42236
rect 71944 42180 72000 42236
rect 72024 42180 72080 42236
rect 72104 42180 72160 42236
rect 71864 42100 71920 42156
rect 71944 42100 72000 42156
rect 72024 42100 72080 42156
rect 72104 42100 72160 42156
rect 71864 42020 71920 42076
rect 71944 42020 72000 42076
rect 72024 42020 72080 42076
rect 72104 42020 72160 42076
rect 71864 41940 71920 41996
rect 71944 41940 72000 41996
rect 72024 41940 72080 41996
rect 72104 41940 72160 41996
rect 71864 32180 71920 32236
rect 71944 32180 72000 32236
rect 72024 32180 72080 32236
rect 72104 32180 72160 32236
rect 71864 32122 71920 32156
rect 71944 32122 72000 32156
rect 72024 32122 72080 32156
rect 72104 32122 72160 32156
rect 71864 32100 71910 32122
rect 71910 32100 71920 32122
rect 71944 32100 71974 32122
rect 71974 32100 71986 32122
rect 71986 32100 72000 32122
rect 72024 32100 72038 32122
rect 72038 32100 72050 32122
rect 72050 32100 72080 32122
rect 72104 32100 72114 32122
rect 72114 32100 72160 32122
rect 71864 32070 71910 32076
rect 71910 32070 71920 32076
rect 71944 32070 71974 32076
rect 71974 32070 71986 32076
rect 71986 32070 72000 32076
rect 72024 32070 72038 32076
rect 72038 32070 72050 32076
rect 72050 32070 72080 32076
rect 72104 32070 72114 32076
rect 72114 32070 72160 32076
rect 71864 32020 71920 32070
rect 71944 32020 72000 32070
rect 72024 32020 72080 32070
rect 72104 32020 72160 32070
rect 71864 31940 71920 31996
rect 71944 31940 72000 31996
rect 72024 31940 72080 31996
rect 72104 31940 72160 31996
rect 71864 22180 71920 22236
rect 71944 22180 72000 22236
rect 72024 22180 72080 22236
rect 72104 22180 72160 22236
rect 71864 22100 71920 22156
rect 71944 22100 72000 22156
rect 72024 22100 72080 22156
rect 72104 22100 72160 22156
rect 71864 22020 71920 22076
rect 71944 22020 72000 22076
rect 72024 22020 72080 22076
rect 72104 22020 72160 22076
rect 71864 21940 71920 21996
rect 71944 21940 72000 21996
rect 72024 21940 72080 21996
rect 72104 21940 72160 21996
rect 71864 12180 71920 12236
rect 71944 12180 72000 12236
rect 72024 12180 72080 12236
rect 72104 12180 72160 12236
rect 71864 12100 71920 12156
rect 71944 12100 72000 12156
rect 72024 12100 72080 12156
rect 72104 12100 72160 12156
rect 71864 12020 71920 12076
rect 71944 12020 72000 12076
rect 72024 12020 72080 12076
rect 72104 12020 72160 12076
rect 71864 11940 71920 11996
rect 71944 11940 72000 11996
rect 72024 11940 72080 11996
rect 72104 11940 72160 11996
rect 74216 84532 74272 84588
rect 74296 84532 74352 84588
rect 74376 84532 74432 84588
rect 74456 84532 74512 84588
rect 74216 84452 74272 84508
rect 74296 84452 74352 84508
rect 74376 84452 74432 84508
rect 74456 84452 74512 84508
rect 74216 84372 74272 84428
rect 74296 84372 74352 84428
rect 74376 84372 74432 84428
rect 74456 84372 74512 84428
rect 74216 84292 74272 84348
rect 74296 84292 74352 84348
rect 74376 84292 74432 84348
rect 74456 84292 74512 84348
rect 74216 74532 74272 74588
rect 74296 74532 74352 74588
rect 74376 74532 74432 74588
rect 74456 74532 74512 74588
rect 74216 74452 74272 74508
rect 74296 74452 74352 74508
rect 74376 74452 74432 74508
rect 74456 74452 74512 74508
rect 74216 74372 74272 74428
rect 74296 74372 74352 74428
rect 74376 74372 74432 74428
rect 74456 74372 74512 74428
rect 74216 74292 74272 74348
rect 74296 74292 74352 74348
rect 74376 74292 74432 74348
rect 74456 74292 74512 74348
rect 74216 64532 74272 64588
rect 74296 64532 74352 64588
rect 74376 64532 74432 64588
rect 74456 64532 74512 64588
rect 74216 64452 74272 64508
rect 74296 64452 74352 64508
rect 74376 64452 74432 64508
rect 74456 64452 74512 64508
rect 74216 64372 74272 64428
rect 74296 64372 74352 64428
rect 74376 64372 74432 64428
rect 74456 64372 74512 64428
rect 74216 64292 74272 64348
rect 74296 64292 74352 64348
rect 74376 64292 74432 64348
rect 74456 64292 74512 64348
rect 74216 54532 74272 54588
rect 74296 54532 74352 54588
rect 74376 54532 74432 54588
rect 74456 54532 74512 54588
rect 74216 54452 74272 54508
rect 74296 54452 74352 54508
rect 74376 54452 74432 54508
rect 74456 54452 74512 54508
rect 74216 54426 74272 54428
rect 74296 54426 74352 54428
rect 74376 54426 74432 54428
rect 74456 54426 74512 54428
rect 74216 54374 74262 54426
rect 74262 54374 74272 54426
rect 74296 54374 74326 54426
rect 74326 54374 74338 54426
rect 74338 54374 74352 54426
rect 74376 54374 74390 54426
rect 74390 54374 74402 54426
rect 74402 54374 74432 54426
rect 74456 54374 74466 54426
rect 74466 54374 74512 54426
rect 74216 54372 74272 54374
rect 74296 54372 74352 54374
rect 74376 54372 74432 54374
rect 74456 54372 74512 54374
rect 74216 54292 74272 54348
rect 74296 54292 74352 54348
rect 74376 54292 74432 54348
rect 74456 54292 74512 54348
rect 74216 44582 74262 44588
rect 74262 44582 74272 44588
rect 74296 44582 74326 44588
rect 74326 44582 74338 44588
rect 74338 44582 74352 44588
rect 74376 44582 74390 44588
rect 74390 44582 74402 44588
rect 74402 44582 74432 44588
rect 74456 44582 74466 44588
rect 74466 44582 74512 44588
rect 74216 44532 74272 44582
rect 74296 44532 74352 44582
rect 74376 44532 74432 44582
rect 74456 44532 74512 44582
rect 74216 44452 74272 44508
rect 74296 44452 74352 44508
rect 74376 44452 74432 44508
rect 74456 44452 74512 44508
rect 74216 44372 74272 44428
rect 74296 44372 74352 44428
rect 74376 44372 74432 44428
rect 74456 44372 74512 44428
rect 74216 44292 74272 44348
rect 74296 44292 74352 44348
rect 74376 44292 74432 44348
rect 74456 44292 74512 44348
rect 74216 34532 74272 34588
rect 74296 34532 74352 34588
rect 74376 34532 74432 34588
rect 74456 34532 74512 34588
rect 74216 34452 74272 34508
rect 74296 34452 74352 34508
rect 74376 34452 74432 34508
rect 74456 34452 74512 34508
rect 74216 34372 74272 34428
rect 74296 34372 74352 34428
rect 74376 34372 74432 34428
rect 74456 34372 74512 34428
rect 74216 34292 74272 34348
rect 74296 34292 74352 34348
rect 74376 34292 74432 34348
rect 74456 34292 74512 34348
rect 74216 24532 74272 24588
rect 74296 24532 74352 24588
rect 74376 24532 74432 24588
rect 74456 24532 74512 24588
rect 74216 24452 74272 24508
rect 74296 24452 74352 24508
rect 74376 24452 74432 24508
rect 74456 24452 74512 24508
rect 74216 24372 74272 24428
rect 74296 24372 74352 24428
rect 74376 24372 74432 24428
rect 74456 24372 74512 24428
rect 74216 24292 74272 24348
rect 74296 24292 74352 24348
rect 74376 24292 74432 24348
rect 74456 24292 74512 24348
rect 74216 14532 74272 14588
rect 74296 14532 74352 14588
rect 74376 14532 74432 14588
rect 74456 14532 74512 14588
rect 74216 14452 74272 14508
rect 74296 14452 74352 14508
rect 74376 14452 74432 14508
rect 74456 14452 74512 14508
rect 74216 14372 74272 14428
rect 74296 14372 74352 14428
rect 74376 14372 74432 14428
rect 74456 14372 74512 14428
rect 74216 14292 74272 14348
rect 74296 14292 74352 14348
rect 74376 14292 74432 14348
rect 74456 14292 74512 14348
rect 74216 4532 74272 4588
rect 74296 4532 74352 4588
rect 74376 4532 74432 4588
rect 74456 4532 74512 4588
rect 74216 4452 74272 4508
rect 74296 4452 74352 4508
rect 74376 4452 74432 4508
rect 74456 4452 74512 4508
rect 74216 4378 74272 4428
rect 74296 4378 74352 4428
rect 74376 4378 74432 4428
rect 74456 4378 74512 4428
rect 74216 4372 74262 4378
rect 74262 4372 74272 4378
rect 74296 4372 74326 4378
rect 74326 4372 74338 4378
rect 74338 4372 74352 4378
rect 74376 4372 74390 4378
rect 74390 4372 74402 4378
rect 74402 4372 74432 4378
rect 74456 4372 74466 4378
rect 74466 4372 74512 4378
rect 74216 4326 74262 4348
rect 74262 4326 74272 4348
rect 74296 4326 74326 4348
rect 74326 4326 74338 4348
rect 74338 4326 74352 4348
rect 74376 4326 74390 4348
rect 74390 4326 74402 4348
rect 74402 4326 74432 4348
rect 74456 4326 74466 4348
rect 74466 4326 74512 4348
rect 74216 4292 74272 4326
rect 74296 4292 74352 4326
rect 74376 4292 74432 4326
rect 74456 4292 74512 4326
rect 71864 2180 71920 2236
rect 71944 2180 72000 2236
rect 72024 2180 72080 2236
rect 72104 2180 72160 2236
rect 71864 2100 71920 2156
rect 71944 2100 72000 2156
rect 72024 2100 72080 2156
rect 72104 2100 72160 2156
rect 71864 2020 71920 2076
rect 71944 2020 72000 2076
rect 72024 2020 72080 2076
rect 72104 2020 72160 2076
rect 71864 1940 71920 1996
rect 71944 1940 72000 1996
rect 72024 1940 72080 1996
rect 72104 1940 72160 1996
<< metal3 >>
rect 964 84592 75028 84616
rect 964 84588 4740 84592
rect 964 84532 2044 84588
rect 2100 84532 4740 84588
rect 964 84528 4740 84532
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84588 10740 84592
rect 5284 84532 5540 84588
rect 5596 84532 8430 84588
rect 8486 84532 10740 84588
rect 5284 84528 10740 84532
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84588 16740 84592
rect 11284 84532 11320 84588
rect 11376 84532 14210 84588
rect 14266 84532 16740 84588
rect 11284 84528 16740 84532
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84588 17140 84592
rect 17124 84528 17140 84532
rect 17204 84528 17220 84592
rect 17284 84588 22740 84592
rect 17284 84532 19990 84588
rect 20046 84532 22740 84588
rect 17284 84528 22740 84532
rect 22804 84528 22820 84592
rect 22884 84588 22900 84592
rect 22884 84528 22900 84532
rect 22964 84528 22980 84592
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84588 28740 84592
rect 23284 84532 25770 84588
rect 25826 84532 28660 84588
rect 28716 84532 28740 84588
rect 23284 84528 28740 84532
rect 28804 84528 28820 84592
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84588 34740 84592
rect 29284 84532 31550 84588
rect 31606 84532 34440 84588
rect 34496 84532 34740 84588
rect 29284 84528 34740 84532
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84588 40740 84592
rect 35284 84532 37330 84588
rect 37386 84532 40220 84588
rect 40276 84532 40740 84588
rect 35284 84528 40740 84532
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84588 46740 84592
rect 41284 84532 43110 84588
rect 43166 84532 46000 84588
rect 46056 84532 46740 84588
rect 41284 84528 46740 84532
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84588 52740 84592
rect 47284 84532 49008 84588
rect 49064 84532 52237 84588
rect 52293 84532 52740 84588
rect 47284 84528 52740 84532
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84588 58740 84592
rect 53284 84532 53638 84588
rect 53694 84532 53806 84588
rect 53862 84532 54550 84588
rect 54606 84532 54940 84588
rect 54996 84532 55656 84588
rect 55712 84532 56234 84588
rect 56290 84532 56679 84588
rect 56735 84532 56983 84588
rect 57039 84532 57825 84588
rect 57881 84532 58465 84588
rect 58521 84532 58740 84588
rect 53284 84528 58740 84532
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84588 59060 84592
rect 59044 84532 59048 84588
rect 59044 84528 59060 84532
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84588 64740 84592
rect 59284 84532 60326 84588
rect 60382 84532 60484 84588
rect 60540 84532 62528 84588
rect 62584 84532 62608 84588
rect 62664 84532 64740 84588
rect 59284 84528 64740 84532
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84588 75028 84592
rect 71284 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 75028 84588
rect 71284 84528 75028 84532
rect 964 84512 75028 84528
rect 964 84508 4740 84512
rect 964 84452 2044 84508
rect 2100 84452 4740 84508
rect 964 84448 4740 84452
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84508 10740 84512
rect 5284 84452 5540 84508
rect 5596 84452 8430 84508
rect 8486 84452 10740 84508
rect 5284 84448 10740 84452
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84508 16740 84512
rect 11284 84452 11320 84508
rect 11376 84452 14210 84508
rect 14266 84452 16740 84508
rect 11284 84448 16740 84452
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84508 17140 84512
rect 17124 84448 17140 84452
rect 17204 84448 17220 84512
rect 17284 84508 22740 84512
rect 17284 84452 19990 84508
rect 20046 84452 22740 84508
rect 17284 84448 22740 84452
rect 22804 84448 22820 84512
rect 22884 84508 22900 84512
rect 22884 84448 22900 84452
rect 22964 84448 22980 84512
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84508 28740 84512
rect 23284 84452 25770 84508
rect 25826 84452 28660 84508
rect 28716 84452 28740 84508
rect 23284 84448 28740 84452
rect 28804 84448 28820 84512
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84508 34740 84512
rect 29284 84452 31550 84508
rect 31606 84452 34440 84508
rect 34496 84452 34740 84508
rect 29284 84448 34740 84452
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84508 40740 84512
rect 35284 84452 37330 84508
rect 37386 84452 40220 84508
rect 40276 84452 40740 84508
rect 35284 84448 40740 84452
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84508 46740 84512
rect 41284 84452 43110 84508
rect 43166 84452 46000 84508
rect 46056 84452 46740 84508
rect 41284 84448 46740 84452
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84508 52740 84512
rect 47284 84452 49008 84508
rect 49064 84452 52237 84508
rect 52293 84452 52740 84508
rect 47284 84448 52740 84452
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84508 58740 84512
rect 53284 84452 53638 84508
rect 53694 84452 53806 84508
rect 53862 84452 54550 84508
rect 54606 84452 54940 84508
rect 54996 84452 55656 84508
rect 55712 84452 56234 84508
rect 56290 84452 56679 84508
rect 56735 84452 56983 84508
rect 57039 84452 57825 84508
rect 57881 84452 58465 84508
rect 58521 84452 58740 84508
rect 53284 84448 58740 84452
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84508 59060 84512
rect 59044 84452 59048 84508
rect 59044 84448 59060 84452
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84508 64740 84512
rect 59284 84452 60326 84508
rect 60382 84452 60484 84508
rect 60540 84452 62528 84508
rect 62584 84452 62608 84508
rect 62664 84452 64740 84508
rect 59284 84448 64740 84452
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84508 75028 84512
rect 71284 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 75028 84508
rect 71284 84448 75028 84452
rect 964 84432 75028 84448
rect 964 84428 4740 84432
rect 964 84372 2044 84428
rect 2100 84372 4740 84428
rect 964 84368 4740 84372
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84428 10740 84432
rect 5284 84372 5540 84428
rect 5596 84372 8430 84428
rect 8486 84372 10740 84428
rect 5284 84368 10740 84372
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84428 16740 84432
rect 11284 84372 11320 84428
rect 11376 84372 14210 84428
rect 14266 84372 16740 84428
rect 11284 84368 16740 84372
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84428 17140 84432
rect 17124 84368 17140 84372
rect 17204 84368 17220 84432
rect 17284 84428 22740 84432
rect 17284 84372 19990 84428
rect 20046 84372 22740 84428
rect 17284 84368 22740 84372
rect 22804 84368 22820 84432
rect 22884 84428 22900 84432
rect 22884 84368 22900 84372
rect 22964 84368 22980 84432
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84428 28740 84432
rect 23284 84372 25770 84428
rect 25826 84372 28660 84428
rect 28716 84372 28740 84428
rect 23284 84368 28740 84372
rect 28804 84368 28820 84432
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84428 34740 84432
rect 29284 84372 31550 84428
rect 31606 84372 34440 84428
rect 34496 84372 34740 84428
rect 29284 84368 34740 84372
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84428 40740 84432
rect 35284 84372 37330 84428
rect 37386 84372 40220 84428
rect 40276 84372 40740 84428
rect 35284 84368 40740 84372
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84428 46740 84432
rect 41284 84372 43110 84428
rect 43166 84372 46000 84428
rect 46056 84372 46740 84428
rect 41284 84368 46740 84372
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84428 52740 84432
rect 47284 84372 49008 84428
rect 49064 84372 52237 84428
rect 52293 84372 52740 84428
rect 47284 84368 52740 84372
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84428 58740 84432
rect 53284 84372 53638 84428
rect 53694 84372 53806 84428
rect 53862 84372 54550 84428
rect 54606 84372 54940 84428
rect 54996 84372 55656 84428
rect 55712 84372 56234 84428
rect 56290 84372 56679 84428
rect 56735 84372 56983 84428
rect 57039 84372 57825 84428
rect 57881 84372 58465 84428
rect 58521 84372 58740 84428
rect 53284 84368 58740 84372
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84428 59060 84432
rect 59044 84372 59048 84428
rect 59044 84368 59060 84372
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84428 64740 84432
rect 59284 84372 60326 84428
rect 60382 84372 60484 84428
rect 60540 84372 62528 84428
rect 62584 84372 62608 84428
rect 62664 84372 64740 84428
rect 59284 84368 64740 84372
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84428 75028 84432
rect 71284 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 75028 84428
rect 71284 84368 75028 84372
rect 964 84352 75028 84368
rect 964 84348 4740 84352
rect 964 84292 2044 84348
rect 2100 84292 4740 84348
rect 964 84288 4740 84292
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84348 10740 84352
rect 5284 84292 5540 84348
rect 5596 84292 8430 84348
rect 8486 84292 10740 84348
rect 5284 84288 10740 84292
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84348 16740 84352
rect 11284 84292 11320 84348
rect 11376 84292 14210 84348
rect 14266 84292 16740 84348
rect 11284 84288 16740 84292
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84348 17140 84352
rect 17124 84288 17140 84292
rect 17204 84288 17220 84352
rect 17284 84348 22740 84352
rect 17284 84292 19990 84348
rect 20046 84292 22740 84348
rect 17284 84288 22740 84292
rect 22804 84288 22820 84352
rect 22884 84348 22900 84352
rect 22884 84288 22900 84292
rect 22964 84288 22980 84352
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84348 28740 84352
rect 23284 84292 25770 84348
rect 25826 84292 28660 84348
rect 28716 84292 28740 84348
rect 23284 84288 28740 84292
rect 28804 84288 28820 84352
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84348 34740 84352
rect 29284 84292 31550 84348
rect 31606 84292 34440 84348
rect 34496 84292 34740 84348
rect 29284 84288 34740 84292
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84348 40740 84352
rect 35284 84292 37330 84348
rect 37386 84292 40220 84348
rect 40276 84292 40740 84348
rect 35284 84288 40740 84292
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84348 46740 84352
rect 41284 84292 43110 84348
rect 43166 84292 46000 84348
rect 46056 84292 46740 84348
rect 41284 84288 46740 84292
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84348 52740 84352
rect 47284 84292 49008 84348
rect 49064 84292 52237 84348
rect 52293 84292 52740 84348
rect 47284 84288 52740 84292
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84348 58740 84352
rect 53284 84292 53638 84348
rect 53694 84292 53806 84348
rect 53862 84292 54550 84348
rect 54606 84292 54940 84348
rect 54996 84292 55656 84348
rect 55712 84292 56234 84348
rect 56290 84292 56679 84348
rect 56735 84292 56983 84348
rect 57039 84292 57825 84348
rect 57881 84292 58465 84348
rect 58521 84292 58740 84348
rect 53284 84288 58740 84292
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84348 59060 84352
rect 59044 84292 59048 84348
rect 59044 84288 59060 84292
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84348 64740 84352
rect 59284 84292 60326 84348
rect 60382 84292 60484 84348
rect 60540 84292 62528 84348
rect 62584 84292 62608 84348
rect 62664 84292 64740 84348
rect 59284 84288 64740 84292
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84348 75028 84352
rect 71284 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 75028 84348
rect 71284 84288 75028 84292
rect 964 84264 75028 84288
rect 964 82240 75028 82264
rect 964 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82236 2220 82240
rect 2284 82236 7740 82240
rect 2320 82180 5393 82236
rect 5449 82180 7740 82236
rect 2204 82176 2220 82180
rect 2284 82176 7740 82180
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82236 13740 82240
rect 8339 82180 11173 82236
rect 11229 82180 13740 82236
rect 8284 82176 13740 82180
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82176 14220 82240
rect 14284 82236 19740 82240
rect 14284 82180 16953 82236
rect 17009 82180 19740 82236
rect 14284 82176 19740 82180
rect 19804 82176 19820 82240
rect 19884 82236 19900 82240
rect 19899 82180 19900 82236
rect 19884 82176 19900 82180
rect 19964 82176 19980 82240
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82236 25740 82240
rect 20284 82180 22733 82236
rect 22789 82180 25623 82236
rect 25679 82180 25740 82236
rect 20284 82176 25740 82180
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82236 31740 82240
rect 26284 82180 28513 82236
rect 28569 82180 31403 82236
rect 31459 82180 31740 82236
rect 26284 82176 31740 82180
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82236 37740 82240
rect 32284 82180 34293 82236
rect 34349 82180 37183 82236
rect 37239 82180 37740 82236
rect 32284 82176 37740 82180
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82236 43740 82240
rect 38284 82180 40073 82236
rect 40129 82180 42963 82236
rect 43019 82180 43740 82236
rect 38284 82176 43740 82180
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82236 49740 82240
rect 44284 82180 45853 82236
rect 45909 82180 48800 82236
rect 48856 82180 49662 82236
rect 49718 82180 49740 82236
rect 44284 82176 49740 82180
rect 49804 82176 49820 82240
rect 49884 82176 49900 82240
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82236 55740 82240
rect 50284 82180 52956 82236
rect 53012 82180 53114 82236
rect 53170 82180 53470 82236
rect 53526 82180 54788 82236
rect 54844 82180 55381 82236
rect 55437 82180 55740 82236
rect 50284 82176 55740 82180
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82236 61740 82240
rect 56284 82180 56527 82236
rect 56583 82180 57963 82236
rect 58019 82180 58043 82236
rect 58099 82180 59206 82236
rect 59262 82180 59364 82236
rect 59420 82180 59672 82236
rect 59728 82180 59818 82236
rect 59874 82180 59954 82236
rect 60010 82180 60034 82236
rect 60090 82180 61740 82236
rect 56284 82176 61740 82180
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82236 67740 82240
rect 62284 82180 62326 82236
rect 62382 82180 62406 82236
rect 62462 82180 67740 82236
rect 62284 82176 67740 82180
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82236 73740 82240
rect 68284 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 73740 82236
rect 68284 82176 73740 82180
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 75028 82240
rect 964 82160 75028 82176
rect 964 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82156 2220 82160
rect 2284 82156 7740 82160
rect 2320 82100 5393 82156
rect 5449 82100 7740 82156
rect 2204 82096 2220 82100
rect 2284 82096 7740 82100
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82156 13740 82160
rect 8339 82100 11173 82156
rect 11229 82100 13740 82156
rect 8284 82096 13740 82100
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82096 14220 82160
rect 14284 82156 19740 82160
rect 14284 82100 16953 82156
rect 17009 82100 19740 82156
rect 14284 82096 19740 82100
rect 19804 82096 19820 82160
rect 19884 82156 19900 82160
rect 19899 82100 19900 82156
rect 19884 82096 19900 82100
rect 19964 82096 19980 82160
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82156 25740 82160
rect 20284 82100 22733 82156
rect 22789 82100 25623 82156
rect 25679 82100 25740 82156
rect 20284 82096 25740 82100
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82156 31740 82160
rect 26284 82100 28513 82156
rect 28569 82100 31403 82156
rect 31459 82100 31740 82156
rect 26284 82096 31740 82100
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82156 37740 82160
rect 32284 82100 34293 82156
rect 34349 82100 37183 82156
rect 37239 82100 37740 82156
rect 32284 82096 37740 82100
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82156 43740 82160
rect 38284 82100 40073 82156
rect 40129 82100 42963 82156
rect 43019 82100 43740 82156
rect 38284 82096 43740 82100
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82156 49740 82160
rect 44284 82100 45853 82156
rect 45909 82100 48800 82156
rect 48856 82100 49662 82156
rect 49718 82100 49740 82156
rect 44284 82096 49740 82100
rect 49804 82096 49820 82160
rect 49884 82096 49900 82160
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82156 55740 82160
rect 50284 82100 52956 82156
rect 53012 82100 53114 82156
rect 53170 82100 53470 82156
rect 53526 82100 54788 82156
rect 54844 82100 55381 82156
rect 55437 82100 55740 82156
rect 50284 82096 55740 82100
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82156 61740 82160
rect 56284 82100 56527 82156
rect 56583 82100 57963 82156
rect 58019 82100 58043 82156
rect 58099 82100 59206 82156
rect 59262 82100 59364 82156
rect 59420 82100 59672 82156
rect 59728 82100 59818 82156
rect 59874 82100 59954 82156
rect 60010 82100 60034 82156
rect 60090 82100 61740 82156
rect 56284 82096 61740 82100
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82156 67740 82160
rect 62284 82100 62326 82156
rect 62382 82100 62406 82156
rect 62462 82100 67740 82156
rect 62284 82096 67740 82100
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82156 73740 82160
rect 68284 82100 71864 82156
rect 71920 82100 71944 82156
rect 72000 82100 72024 82156
rect 72080 82100 72104 82156
rect 72160 82100 73740 82156
rect 68284 82096 73740 82100
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 75028 82160
rect 964 82080 75028 82096
rect 964 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82076 2220 82080
rect 2284 82076 7740 82080
rect 2320 82020 5393 82076
rect 5449 82020 7740 82076
rect 2204 82016 2220 82020
rect 2284 82016 7740 82020
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82076 13740 82080
rect 8339 82020 11173 82076
rect 11229 82020 13740 82076
rect 8284 82016 13740 82020
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82016 14220 82080
rect 14284 82076 19740 82080
rect 14284 82020 16953 82076
rect 17009 82020 19740 82076
rect 14284 82016 19740 82020
rect 19804 82016 19820 82080
rect 19884 82076 19900 82080
rect 19899 82020 19900 82076
rect 19884 82016 19900 82020
rect 19964 82016 19980 82080
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82076 25740 82080
rect 20284 82020 22733 82076
rect 22789 82020 25623 82076
rect 25679 82020 25740 82076
rect 20284 82016 25740 82020
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82076 31740 82080
rect 26284 82020 28513 82076
rect 28569 82020 31403 82076
rect 31459 82020 31740 82076
rect 26284 82016 31740 82020
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82076 37740 82080
rect 32284 82020 34293 82076
rect 34349 82020 37183 82076
rect 37239 82020 37740 82076
rect 32284 82016 37740 82020
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82076 43740 82080
rect 38284 82020 40073 82076
rect 40129 82020 42963 82076
rect 43019 82020 43740 82076
rect 38284 82016 43740 82020
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82076 49740 82080
rect 44284 82020 45853 82076
rect 45909 82020 48800 82076
rect 48856 82020 49662 82076
rect 49718 82020 49740 82076
rect 44284 82016 49740 82020
rect 49804 82016 49820 82080
rect 49884 82016 49900 82080
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82076 55740 82080
rect 50284 82020 52956 82076
rect 53012 82020 53114 82076
rect 53170 82020 53470 82076
rect 53526 82020 54788 82076
rect 54844 82020 55381 82076
rect 55437 82020 55740 82076
rect 50284 82016 55740 82020
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82076 61740 82080
rect 56284 82020 56527 82076
rect 56583 82020 57963 82076
rect 58019 82020 58043 82076
rect 58099 82020 59206 82076
rect 59262 82020 59364 82076
rect 59420 82020 59672 82076
rect 59728 82020 59818 82076
rect 59874 82020 59954 82076
rect 60010 82020 60034 82076
rect 60090 82020 61740 82076
rect 56284 82016 61740 82020
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82076 67740 82080
rect 62284 82020 62326 82076
rect 62382 82020 62406 82076
rect 62462 82020 67740 82076
rect 62284 82016 67740 82020
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82076 73740 82080
rect 68284 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 73740 82076
rect 68284 82016 73740 82020
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 75028 82080
rect 964 82000 75028 82016
rect 964 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81996 2220 82000
rect 2284 81996 7740 82000
rect 2320 81940 5393 81996
rect 5449 81940 7740 81996
rect 2204 81936 2220 81940
rect 2284 81936 7740 81940
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81996 13740 82000
rect 8339 81940 11173 81996
rect 11229 81940 13740 81996
rect 8284 81936 13740 81940
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81936 14220 82000
rect 14284 81996 19740 82000
rect 14284 81940 16953 81996
rect 17009 81940 19740 81996
rect 14284 81936 19740 81940
rect 19804 81936 19820 82000
rect 19884 81996 19900 82000
rect 19899 81940 19900 81996
rect 19884 81936 19900 81940
rect 19964 81936 19980 82000
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81996 25740 82000
rect 20284 81940 22733 81996
rect 22789 81940 25623 81996
rect 25679 81940 25740 81996
rect 20284 81936 25740 81940
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81996 31740 82000
rect 26284 81940 28513 81996
rect 28569 81940 31403 81996
rect 31459 81940 31740 81996
rect 26284 81936 31740 81940
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81996 37740 82000
rect 32284 81940 34293 81996
rect 34349 81940 37183 81996
rect 37239 81940 37740 81996
rect 32284 81936 37740 81940
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81996 43740 82000
rect 38284 81940 40073 81996
rect 40129 81940 42963 81996
rect 43019 81940 43740 81996
rect 38284 81936 43740 81940
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81996 49740 82000
rect 44284 81940 45853 81996
rect 45909 81940 48800 81996
rect 48856 81940 49662 81996
rect 49718 81940 49740 81996
rect 44284 81936 49740 81940
rect 49804 81936 49820 82000
rect 49884 81936 49900 82000
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81996 55740 82000
rect 50284 81940 52956 81996
rect 53012 81940 53114 81996
rect 53170 81940 53470 81996
rect 53526 81940 54788 81996
rect 54844 81940 55381 81996
rect 55437 81940 55740 81996
rect 50284 81936 55740 81940
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81996 61740 82000
rect 56284 81940 56527 81996
rect 56583 81940 57963 81996
rect 58019 81940 58043 81996
rect 58099 81940 59206 81996
rect 59262 81940 59364 81996
rect 59420 81940 59672 81996
rect 59728 81940 59818 81996
rect 59874 81940 59954 81996
rect 60010 81940 60034 81996
rect 60090 81940 61740 81996
rect 56284 81936 61740 81940
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81996 67740 82000
rect 62284 81940 62326 81996
rect 62382 81940 62406 81996
rect 62462 81940 67740 81996
rect 62284 81936 67740 81940
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81996 73740 82000
rect 68284 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 73740 81996
rect 68284 81936 73740 81940
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 75028 82000
rect 964 81912 75028 81936
rect 964 74592 75028 74616
rect 964 74588 4740 74592
rect 964 74532 2044 74588
rect 2100 74532 4740 74588
rect 964 74528 4740 74532
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74588 10740 74592
rect 5284 74532 5540 74588
rect 5596 74532 8430 74588
rect 8486 74532 10740 74588
rect 5284 74528 10740 74532
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74588 16740 74592
rect 11284 74532 11320 74588
rect 11376 74532 14210 74588
rect 14266 74532 16740 74588
rect 11284 74528 16740 74532
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74588 17140 74592
rect 17124 74528 17140 74532
rect 17204 74528 17220 74592
rect 17284 74588 22740 74592
rect 17284 74532 19990 74588
rect 20046 74532 22740 74588
rect 17284 74528 22740 74532
rect 22804 74528 22820 74592
rect 22884 74588 22900 74592
rect 22884 74528 22900 74532
rect 22964 74528 22980 74592
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74588 28740 74592
rect 23284 74532 25770 74588
rect 25826 74532 28660 74588
rect 28716 74532 28740 74588
rect 23284 74528 28740 74532
rect 28804 74528 28820 74592
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74588 34740 74592
rect 29284 74532 31550 74588
rect 31606 74532 34440 74588
rect 34496 74532 34740 74588
rect 29284 74528 34740 74532
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74588 40740 74592
rect 35284 74532 37330 74588
rect 37386 74532 40220 74588
rect 40276 74532 40740 74588
rect 35284 74528 40740 74532
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74588 46740 74592
rect 41284 74532 43110 74588
rect 43166 74532 46000 74588
rect 46056 74532 46740 74588
rect 41284 74528 46740 74532
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74588 52740 74592
rect 47284 74532 49008 74588
rect 49064 74532 52237 74588
rect 52293 74532 52740 74588
rect 47284 74528 52740 74532
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74588 58740 74592
rect 53284 74532 53638 74588
rect 53694 74532 53806 74588
rect 53862 74532 54550 74588
rect 54606 74532 54940 74588
rect 54996 74532 55656 74588
rect 55712 74532 56234 74588
rect 56290 74532 56679 74588
rect 56735 74532 56983 74588
rect 57039 74532 57825 74588
rect 57881 74532 58465 74588
rect 58521 74532 58740 74588
rect 53284 74528 58740 74532
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74588 59060 74592
rect 59044 74532 59048 74588
rect 59044 74528 59060 74532
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74588 64740 74592
rect 59284 74532 60326 74588
rect 60382 74532 60484 74588
rect 60540 74532 62528 74588
rect 62584 74532 62608 74588
rect 62664 74532 64740 74588
rect 59284 74528 64740 74532
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74588 75028 74592
rect 71284 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 75028 74588
rect 71284 74528 75028 74532
rect 964 74512 75028 74528
rect 964 74508 4740 74512
rect 964 74452 2044 74508
rect 2100 74452 4740 74508
rect 964 74448 4740 74452
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74508 10740 74512
rect 5284 74452 5540 74508
rect 5596 74452 8430 74508
rect 8486 74452 10740 74508
rect 5284 74448 10740 74452
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74508 16740 74512
rect 11284 74452 11320 74508
rect 11376 74452 14210 74508
rect 14266 74452 16740 74508
rect 11284 74448 16740 74452
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74508 17140 74512
rect 17124 74448 17140 74452
rect 17204 74448 17220 74512
rect 17284 74508 22740 74512
rect 17284 74452 19990 74508
rect 20046 74452 22740 74508
rect 17284 74448 22740 74452
rect 22804 74448 22820 74512
rect 22884 74508 22900 74512
rect 22884 74448 22900 74452
rect 22964 74448 22980 74512
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74508 28740 74512
rect 23284 74452 25770 74508
rect 25826 74452 28660 74508
rect 28716 74452 28740 74508
rect 23284 74448 28740 74452
rect 28804 74448 28820 74512
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74508 34740 74512
rect 29284 74452 31550 74508
rect 31606 74452 34440 74508
rect 34496 74452 34740 74508
rect 29284 74448 34740 74452
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74508 40740 74512
rect 35284 74452 37330 74508
rect 37386 74452 40220 74508
rect 40276 74452 40740 74508
rect 35284 74448 40740 74452
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74508 46740 74512
rect 41284 74452 43110 74508
rect 43166 74452 46000 74508
rect 46056 74452 46740 74508
rect 41284 74448 46740 74452
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74508 52740 74512
rect 47284 74452 49008 74508
rect 49064 74452 52237 74508
rect 52293 74452 52740 74508
rect 47284 74448 52740 74452
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74508 58740 74512
rect 53284 74452 53638 74508
rect 53694 74452 53806 74508
rect 53862 74452 54550 74508
rect 54606 74452 54940 74508
rect 54996 74452 55656 74508
rect 55712 74452 56234 74508
rect 56290 74452 56679 74508
rect 56735 74452 56983 74508
rect 57039 74452 57825 74508
rect 57881 74452 58465 74508
rect 58521 74452 58740 74508
rect 53284 74448 58740 74452
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74508 59060 74512
rect 59044 74452 59048 74508
rect 59044 74448 59060 74452
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74508 64740 74512
rect 59284 74452 60326 74508
rect 60382 74452 60484 74508
rect 60540 74452 62528 74508
rect 62584 74452 62608 74508
rect 62664 74452 64740 74508
rect 59284 74448 64740 74452
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74508 75028 74512
rect 71284 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 75028 74508
rect 71284 74448 75028 74452
rect 964 74432 75028 74448
rect 964 74428 4740 74432
rect 964 74372 2044 74428
rect 2100 74372 4740 74428
rect 964 74368 4740 74372
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74428 10740 74432
rect 5284 74372 5540 74428
rect 5596 74372 8430 74428
rect 8486 74372 10740 74428
rect 5284 74368 10740 74372
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74428 16740 74432
rect 11284 74372 11320 74428
rect 11376 74372 14210 74428
rect 14266 74372 16740 74428
rect 11284 74368 16740 74372
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74428 17140 74432
rect 17124 74368 17140 74372
rect 17204 74368 17220 74432
rect 17284 74428 22740 74432
rect 17284 74372 19990 74428
rect 20046 74372 22740 74428
rect 17284 74368 22740 74372
rect 22804 74368 22820 74432
rect 22884 74428 22900 74432
rect 22884 74368 22900 74372
rect 22964 74368 22980 74432
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74428 28740 74432
rect 23284 74372 25770 74428
rect 25826 74372 28660 74428
rect 28716 74372 28740 74428
rect 23284 74368 28740 74372
rect 28804 74368 28820 74432
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74428 34740 74432
rect 29284 74372 31550 74428
rect 31606 74372 34440 74428
rect 34496 74372 34740 74428
rect 29284 74368 34740 74372
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74428 40740 74432
rect 35284 74372 37330 74428
rect 37386 74372 40220 74428
rect 40276 74372 40740 74428
rect 35284 74368 40740 74372
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74428 46740 74432
rect 41284 74372 43110 74428
rect 43166 74372 46000 74428
rect 46056 74372 46740 74428
rect 41284 74368 46740 74372
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74428 52740 74432
rect 47284 74372 49008 74428
rect 49064 74372 52237 74428
rect 52293 74372 52740 74428
rect 47284 74368 52740 74372
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74428 58740 74432
rect 53284 74372 53638 74428
rect 53694 74372 53806 74428
rect 53862 74372 54550 74428
rect 54606 74372 54940 74428
rect 54996 74372 55656 74428
rect 55712 74372 56234 74428
rect 56290 74372 56679 74428
rect 56735 74372 56983 74428
rect 57039 74372 57825 74428
rect 57881 74372 58465 74428
rect 58521 74372 58740 74428
rect 53284 74368 58740 74372
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74428 59060 74432
rect 59044 74372 59048 74428
rect 59044 74368 59060 74372
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74428 64740 74432
rect 59284 74372 60326 74428
rect 60382 74372 60484 74428
rect 60540 74372 62528 74428
rect 62584 74372 62608 74428
rect 62664 74372 64740 74428
rect 59284 74368 64740 74372
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74428 75028 74432
rect 71284 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 75028 74428
rect 71284 74368 75028 74372
rect 964 74352 75028 74368
rect 964 74348 4740 74352
rect 964 74292 2044 74348
rect 2100 74292 4740 74348
rect 964 74288 4740 74292
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74348 10740 74352
rect 5284 74292 5540 74348
rect 5596 74292 8430 74348
rect 8486 74292 10740 74348
rect 5284 74288 10740 74292
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74348 16740 74352
rect 11284 74292 11320 74348
rect 11376 74292 14210 74348
rect 14266 74292 16740 74348
rect 11284 74288 16740 74292
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74348 17140 74352
rect 17124 74288 17140 74292
rect 17204 74288 17220 74352
rect 17284 74348 22740 74352
rect 17284 74292 19990 74348
rect 20046 74292 22740 74348
rect 17284 74288 22740 74292
rect 22804 74288 22820 74352
rect 22884 74348 22900 74352
rect 22884 74288 22900 74292
rect 22964 74288 22980 74352
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74348 28740 74352
rect 23284 74292 25770 74348
rect 25826 74292 28660 74348
rect 28716 74292 28740 74348
rect 23284 74288 28740 74292
rect 28804 74288 28820 74352
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74348 34740 74352
rect 29284 74292 31550 74348
rect 31606 74292 34440 74348
rect 34496 74292 34740 74348
rect 29284 74288 34740 74292
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74348 40740 74352
rect 35284 74292 37330 74348
rect 37386 74292 40220 74348
rect 40276 74292 40740 74348
rect 35284 74288 40740 74292
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74348 46740 74352
rect 41284 74292 43110 74348
rect 43166 74292 46000 74348
rect 46056 74292 46740 74348
rect 41284 74288 46740 74292
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74348 52740 74352
rect 47284 74292 49008 74348
rect 49064 74292 52237 74348
rect 52293 74292 52740 74348
rect 47284 74288 52740 74292
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74348 58740 74352
rect 53284 74292 53638 74348
rect 53694 74292 53806 74348
rect 53862 74292 54550 74348
rect 54606 74292 54940 74348
rect 54996 74292 55656 74348
rect 55712 74292 56234 74348
rect 56290 74292 56679 74348
rect 56735 74292 56983 74348
rect 57039 74292 57825 74348
rect 57881 74292 58465 74348
rect 58521 74292 58740 74348
rect 53284 74288 58740 74292
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74348 59060 74352
rect 59044 74292 59048 74348
rect 59044 74288 59060 74292
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74348 64740 74352
rect 59284 74292 60326 74348
rect 60382 74292 60484 74348
rect 60540 74292 62528 74348
rect 62584 74292 62608 74348
rect 62664 74292 64740 74348
rect 59284 74288 64740 74292
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74348 75028 74352
rect 71284 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 75028 74348
rect 71284 74288 75028 74292
rect 964 74264 75028 74288
rect 964 72240 75028 72264
rect 964 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72236 2220 72240
rect 2284 72236 7740 72240
rect 2320 72180 5393 72236
rect 5449 72180 7740 72236
rect 2204 72176 2220 72180
rect 2284 72176 7740 72180
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72236 13740 72240
rect 8339 72180 11173 72236
rect 11229 72180 13740 72236
rect 8284 72176 13740 72180
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72176 14220 72240
rect 14284 72236 19740 72240
rect 14284 72180 16953 72236
rect 17009 72180 19740 72236
rect 14284 72176 19740 72180
rect 19804 72176 19820 72240
rect 19884 72236 19900 72240
rect 19899 72180 19900 72236
rect 19884 72176 19900 72180
rect 19964 72176 19980 72240
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72236 25740 72240
rect 20284 72180 22733 72236
rect 22789 72180 25623 72236
rect 25679 72180 25740 72236
rect 20284 72176 25740 72180
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72236 31740 72240
rect 26284 72180 28513 72236
rect 28569 72180 31403 72236
rect 31459 72180 31740 72236
rect 26284 72176 31740 72180
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72236 37740 72240
rect 32284 72180 34293 72236
rect 34349 72180 37183 72236
rect 37239 72180 37740 72236
rect 32284 72176 37740 72180
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72236 43740 72240
rect 38284 72180 40073 72236
rect 40129 72180 42963 72236
rect 43019 72180 43740 72236
rect 38284 72176 43740 72180
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72236 49740 72240
rect 44284 72180 45853 72236
rect 45909 72180 48800 72236
rect 48856 72180 49662 72236
rect 49718 72180 49740 72236
rect 44284 72176 49740 72180
rect 49804 72176 49820 72240
rect 49884 72176 49900 72240
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72236 55740 72240
rect 50284 72180 52956 72236
rect 53012 72180 53114 72236
rect 53170 72180 53470 72236
rect 53526 72180 54788 72236
rect 54844 72180 55381 72236
rect 55437 72180 55740 72236
rect 50284 72176 55740 72180
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72236 61740 72240
rect 56284 72180 56527 72236
rect 56583 72180 57963 72236
rect 58019 72180 58043 72236
rect 58099 72180 59206 72236
rect 59262 72180 59364 72236
rect 59420 72180 59672 72236
rect 59728 72180 59818 72236
rect 59874 72180 59954 72236
rect 60010 72180 60034 72236
rect 60090 72180 61740 72236
rect 56284 72176 61740 72180
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72236 67740 72240
rect 62284 72180 62326 72236
rect 62382 72180 62406 72236
rect 62462 72180 67740 72236
rect 62284 72176 67740 72180
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72236 73740 72240
rect 68284 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 73740 72236
rect 68284 72176 73740 72180
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 75028 72240
rect 964 72160 75028 72176
rect 964 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72156 2220 72160
rect 2284 72156 7740 72160
rect 2320 72100 5393 72156
rect 5449 72100 7740 72156
rect 2204 72096 2220 72100
rect 2284 72096 7740 72100
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72156 13740 72160
rect 8339 72100 11173 72156
rect 11229 72100 13740 72156
rect 8284 72096 13740 72100
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72096 14220 72160
rect 14284 72156 19740 72160
rect 14284 72100 16953 72156
rect 17009 72100 19740 72156
rect 14284 72096 19740 72100
rect 19804 72096 19820 72160
rect 19884 72156 19900 72160
rect 19899 72100 19900 72156
rect 19884 72096 19900 72100
rect 19964 72096 19980 72160
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72156 25740 72160
rect 20284 72100 22733 72156
rect 22789 72100 25623 72156
rect 25679 72100 25740 72156
rect 20284 72096 25740 72100
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72156 31740 72160
rect 26284 72100 28513 72156
rect 28569 72100 31403 72156
rect 31459 72100 31740 72156
rect 26284 72096 31740 72100
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72156 37740 72160
rect 32284 72100 34293 72156
rect 34349 72100 37183 72156
rect 37239 72100 37740 72156
rect 32284 72096 37740 72100
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72156 43740 72160
rect 38284 72100 40073 72156
rect 40129 72100 42963 72156
rect 43019 72100 43740 72156
rect 38284 72096 43740 72100
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72156 49740 72160
rect 44284 72100 45853 72156
rect 45909 72100 48800 72156
rect 48856 72100 49662 72156
rect 49718 72100 49740 72156
rect 44284 72096 49740 72100
rect 49804 72096 49820 72160
rect 49884 72096 49900 72160
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72156 55740 72160
rect 50284 72100 52956 72156
rect 53012 72100 53114 72156
rect 53170 72100 53470 72156
rect 53526 72100 54788 72156
rect 54844 72100 55381 72156
rect 55437 72100 55740 72156
rect 50284 72096 55740 72100
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72156 61740 72160
rect 56284 72100 56527 72156
rect 56583 72100 57963 72156
rect 58019 72100 58043 72156
rect 58099 72100 59206 72156
rect 59262 72100 59364 72156
rect 59420 72100 59672 72156
rect 59728 72100 59818 72156
rect 59874 72100 59954 72156
rect 60010 72100 60034 72156
rect 60090 72100 61740 72156
rect 56284 72096 61740 72100
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72156 67740 72160
rect 62284 72100 62326 72156
rect 62382 72100 62406 72156
rect 62462 72100 67740 72156
rect 62284 72096 67740 72100
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72156 73740 72160
rect 68284 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 73740 72156
rect 68284 72096 73740 72100
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 75028 72160
rect 964 72080 75028 72096
rect 964 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72076 2220 72080
rect 2284 72076 7740 72080
rect 2320 72020 5393 72076
rect 5449 72020 7740 72076
rect 2204 72016 2220 72020
rect 2284 72016 7740 72020
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72076 13740 72080
rect 8339 72020 11173 72076
rect 11229 72020 13740 72076
rect 8284 72016 13740 72020
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72016 14220 72080
rect 14284 72076 19740 72080
rect 14284 72020 16953 72076
rect 17009 72020 19740 72076
rect 14284 72016 19740 72020
rect 19804 72016 19820 72080
rect 19884 72076 19900 72080
rect 19899 72020 19900 72076
rect 19884 72016 19900 72020
rect 19964 72016 19980 72080
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72076 25740 72080
rect 20284 72020 22733 72076
rect 22789 72020 25623 72076
rect 25679 72020 25740 72076
rect 20284 72016 25740 72020
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72076 31740 72080
rect 26284 72020 28513 72076
rect 28569 72020 31403 72076
rect 31459 72020 31740 72076
rect 26284 72016 31740 72020
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72076 37740 72080
rect 32284 72020 34293 72076
rect 34349 72020 37183 72076
rect 37239 72020 37740 72076
rect 32284 72016 37740 72020
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72076 43740 72080
rect 38284 72020 40073 72076
rect 40129 72020 42963 72076
rect 43019 72020 43740 72076
rect 38284 72016 43740 72020
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72076 49740 72080
rect 44284 72020 45853 72076
rect 45909 72020 48800 72076
rect 48856 72020 49662 72076
rect 49718 72020 49740 72076
rect 44284 72016 49740 72020
rect 49804 72016 49820 72080
rect 49884 72016 49900 72080
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72076 55740 72080
rect 50284 72020 52956 72076
rect 53012 72020 53114 72076
rect 53170 72020 53470 72076
rect 53526 72020 54788 72076
rect 54844 72020 55381 72076
rect 55437 72020 55740 72076
rect 50284 72016 55740 72020
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72076 61740 72080
rect 56284 72020 56527 72076
rect 56583 72020 57963 72076
rect 58019 72020 58043 72076
rect 58099 72020 59206 72076
rect 59262 72020 59364 72076
rect 59420 72020 59672 72076
rect 59728 72020 59818 72076
rect 59874 72020 59954 72076
rect 60010 72020 60034 72076
rect 60090 72020 61740 72076
rect 56284 72016 61740 72020
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72076 67740 72080
rect 62284 72020 62326 72076
rect 62382 72020 62406 72076
rect 62462 72020 67740 72076
rect 62284 72016 67740 72020
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72076 73740 72080
rect 68284 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 73740 72076
rect 68284 72016 73740 72020
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 75028 72080
rect 964 72000 75028 72016
rect 964 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71996 2220 72000
rect 2284 71996 7740 72000
rect 2320 71940 5393 71996
rect 5449 71940 7740 71996
rect 2204 71936 2220 71940
rect 2284 71936 7740 71940
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71996 13740 72000
rect 8339 71940 11173 71996
rect 11229 71940 13740 71996
rect 8284 71936 13740 71940
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71936 14220 72000
rect 14284 71996 19740 72000
rect 14284 71940 16953 71996
rect 17009 71940 19740 71996
rect 14284 71936 19740 71940
rect 19804 71936 19820 72000
rect 19884 71996 19900 72000
rect 19899 71940 19900 71996
rect 19884 71936 19900 71940
rect 19964 71936 19980 72000
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71996 25740 72000
rect 20284 71940 22733 71996
rect 22789 71940 25623 71996
rect 25679 71940 25740 71996
rect 20284 71936 25740 71940
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71996 31740 72000
rect 26284 71940 28513 71996
rect 28569 71940 31403 71996
rect 31459 71940 31740 71996
rect 26284 71936 31740 71940
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71996 37740 72000
rect 32284 71940 34293 71996
rect 34349 71940 37183 71996
rect 37239 71940 37740 71996
rect 32284 71936 37740 71940
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71996 43740 72000
rect 38284 71940 40073 71996
rect 40129 71940 42963 71996
rect 43019 71940 43740 71996
rect 38284 71936 43740 71940
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71996 49740 72000
rect 44284 71940 45853 71996
rect 45909 71940 48800 71996
rect 48856 71940 49662 71996
rect 49718 71940 49740 71996
rect 44284 71936 49740 71940
rect 49804 71936 49820 72000
rect 49884 71936 49900 72000
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71996 55740 72000
rect 50284 71940 52956 71996
rect 53012 71940 53114 71996
rect 53170 71940 53470 71996
rect 53526 71940 54788 71996
rect 54844 71940 55381 71996
rect 55437 71940 55740 71996
rect 50284 71936 55740 71940
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71996 61740 72000
rect 56284 71940 56527 71996
rect 56583 71940 57963 71996
rect 58019 71940 58043 71996
rect 58099 71940 59206 71996
rect 59262 71940 59364 71996
rect 59420 71940 59672 71996
rect 59728 71940 59818 71996
rect 59874 71940 59954 71996
rect 60010 71940 60034 71996
rect 60090 71940 61740 71996
rect 56284 71936 61740 71940
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71996 67740 72000
rect 62284 71940 62326 71996
rect 62382 71940 62406 71996
rect 62462 71940 67740 71996
rect 62284 71936 67740 71940
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71996 73740 72000
rect 68284 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 73740 71996
rect 68284 71936 73740 71940
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 75028 72000
rect 964 71912 75028 71936
rect 964 64592 75028 64616
rect 964 64588 4740 64592
rect 964 64532 2044 64588
rect 2100 64532 4740 64588
rect 964 64528 4740 64532
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64588 10740 64592
rect 5284 64532 5540 64588
rect 5596 64532 8430 64588
rect 8486 64532 10740 64588
rect 5284 64528 10740 64532
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64588 16740 64592
rect 11284 64532 11320 64588
rect 11376 64532 14210 64588
rect 14266 64532 16740 64588
rect 11284 64528 16740 64532
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64588 17140 64592
rect 17124 64528 17140 64532
rect 17204 64528 17220 64592
rect 17284 64588 22740 64592
rect 17284 64532 19990 64588
rect 20046 64532 22740 64588
rect 17284 64528 22740 64532
rect 22804 64528 22820 64592
rect 22884 64588 22900 64592
rect 22884 64528 22900 64532
rect 22964 64528 22980 64592
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64588 28740 64592
rect 23284 64532 25770 64588
rect 25826 64532 28660 64588
rect 28716 64532 28740 64588
rect 23284 64528 28740 64532
rect 28804 64528 28820 64592
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64588 34740 64592
rect 29284 64532 31550 64588
rect 31606 64532 34440 64588
rect 34496 64532 34740 64588
rect 29284 64528 34740 64532
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64588 40740 64592
rect 35284 64532 37330 64588
rect 37386 64532 40220 64588
rect 40276 64532 40740 64588
rect 35284 64528 40740 64532
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64588 46740 64592
rect 41284 64532 43110 64588
rect 43166 64532 46000 64588
rect 46056 64532 46740 64588
rect 41284 64528 46740 64532
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64588 52740 64592
rect 47284 64532 49008 64588
rect 49064 64532 52237 64588
rect 52293 64532 52740 64588
rect 47284 64528 52740 64532
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64588 58740 64592
rect 53284 64532 53638 64588
rect 53694 64532 53806 64588
rect 53862 64532 54550 64588
rect 54606 64532 54940 64588
rect 54996 64532 55656 64588
rect 55712 64532 56234 64588
rect 56290 64532 56679 64588
rect 56735 64532 56983 64588
rect 57039 64532 57825 64588
rect 57881 64532 58465 64588
rect 58521 64532 58740 64588
rect 53284 64528 58740 64532
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64588 59060 64592
rect 59044 64532 59048 64588
rect 59044 64528 59060 64532
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64588 64740 64592
rect 59284 64532 60326 64588
rect 60382 64532 60484 64588
rect 60540 64532 62528 64588
rect 62584 64532 62608 64588
rect 62664 64532 64740 64588
rect 59284 64528 64740 64532
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64588 75028 64592
rect 71284 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 75028 64588
rect 71284 64528 75028 64532
rect 964 64512 75028 64528
rect 964 64508 4740 64512
rect 964 64452 2044 64508
rect 2100 64452 4740 64508
rect 964 64448 4740 64452
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64508 10740 64512
rect 5284 64452 5540 64508
rect 5596 64452 8430 64508
rect 8486 64452 10740 64508
rect 5284 64448 10740 64452
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64508 16740 64512
rect 11284 64452 11320 64508
rect 11376 64452 14210 64508
rect 14266 64452 16740 64508
rect 11284 64448 16740 64452
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64508 17140 64512
rect 17124 64448 17140 64452
rect 17204 64448 17220 64512
rect 17284 64508 22740 64512
rect 17284 64452 19990 64508
rect 20046 64452 22740 64508
rect 17284 64448 22740 64452
rect 22804 64448 22820 64512
rect 22884 64508 22900 64512
rect 22884 64448 22900 64452
rect 22964 64448 22980 64512
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64508 28740 64512
rect 23284 64452 25770 64508
rect 25826 64452 28660 64508
rect 28716 64452 28740 64508
rect 23284 64448 28740 64452
rect 28804 64448 28820 64512
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64508 34740 64512
rect 29284 64452 31550 64508
rect 31606 64452 34440 64508
rect 34496 64452 34740 64508
rect 29284 64448 34740 64452
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64508 40740 64512
rect 35284 64452 37330 64508
rect 37386 64452 40220 64508
rect 40276 64452 40740 64508
rect 35284 64448 40740 64452
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64508 46740 64512
rect 41284 64452 43110 64508
rect 43166 64452 46000 64508
rect 46056 64452 46740 64508
rect 41284 64448 46740 64452
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64508 52740 64512
rect 47284 64452 49008 64508
rect 49064 64452 52237 64508
rect 52293 64452 52740 64508
rect 47284 64448 52740 64452
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64508 58740 64512
rect 53284 64452 53638 64508
rect 53694 64452 53806 64508
rect 53862 64452 54550 64508
rect 54606 64452 54940 64508
rect 54996 64452 55656 64508
rect 55712 64452 56234 64508
rect 56290 64452 56679 64508
rect 56735 64452 56983 64508
rect 57039 64452 57825 64508
rect 57881 64452 58465 64508
rect 58521 64452 58740 64508
rect 53284 64448 58740 64452
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64508 59060 64512
rect 59044 64452 59048 64508
rect 59044 64448 59060 64452
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64508 64740 64512
rect 59284 64452 60326 64508
rect 60382 64452 60484 64508
rect 60540 64452 62528 64508
rect 62584 64452 62608 64508
rect 62664 64452 64740 64508
rect 59284 64448 64740 64452
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64508 75028 64512
rect 71284 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 75028 64508
rect 71284 64448 75028 64452
rect 964 64432 75028 64448
rect 964 64428 4740 64432
rect 964 64372 2044 64428
rect 2100 64372 4740 64428
rect 964 64368 4740 64372
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64428 10740 64432
rect 5284 64372 5540 64428
rect 5596 64372 8430 64428
rect 8486 64372 10740 64428
rect 5284 64368 10740 64372
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64428 16740 64432
rect 11284 64372 11320 64428
rect 11376 64372 14210 64428
rect 14266 64372 16740 64428
rect 11284 64368 16740 64372
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64428 17140 64432
rect 17124 64368 17140 64372
rect 17204 64368 17220 64432
rect 17284 64428 22740 64432
rect 17284 64372 19990 64428
rect 20046 64372 22740 64428
rect 17284 64368 22740 64372
rect 22804 64368 22820 64432
rect 22884 64428 22900 64432
rect 22884 64368 22900 64372
rect 22964 64368 22980 64432
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64428 28740 64432
rect 23284 64372 25770 64428
rect 25826 64372 28660 64428
rect 28716 64372 28740 64428
rect 23284 64368 28740 64372
rect 28804 64368 28820 64432
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64428 34740 64432
rect 29284 64372 31550 64428
rect 31606 64372 34440 64428
rect 34496 64372 34740 64428
rect 29284 64368 34740 64372
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64428 40740 64432
rect 35284 64372 37330 64428
rect 37386 64372 40220 64428
rect 40276 64372 40740 64428
rect 35284 64368 40740 64372
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64428 46740 64432
rect 41284 64372 43110 64428
rect 43166 64372 46000 64428
rect 46056 64372 46740 64428
rect 41284 64368 46740 64372
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64428 52740 64432
rect 47284 64372 49008 64428
rect 49064 64372 52237 64428
rect 52293 64372 52740 64428
rect 47284 64368 52740 64372
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64428 58740 64432
rect 53284 64372 53638 64428
rect 53694 64372 53806 64428
rect 53862 64372 54550 64428
rect 54606 64372 54940 64428
rect 54996 64372 55656 64428
rect 55712 64372 56234 64428
rect 56290 64372 56679 64428
rect 56735 64372 56983 64428
rect 57039 64372 57825 64428
rect 57881 64372 58465 64428
rect 58521 64372 58740 64428
rect 53284 64368 58740 64372
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64428 59060 64432
rect 59044 64372 59048 64428
rect 59044 64368 59060 64372
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64428 64740 64432
rect 59284 64372 60326 64428
rect 60382 64372 60484 64428
rect 60540 64372 62528 64428
rect 62584 64372 62608 64428
rect 62664 64372 64740 64428
rect 59284 64368 64740 64372
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64428 75028 64432
rect 71284 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 75028 64428
rect 71284 64368 75028 64372
rect 964 64352 75028 64368
rect 964 64348 4740 64352
rect 964 64292 2044 64348
rect 2100 64292 4740 64348
rect 964 64288 4740 64292
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64348 10740 64352
rect 5284 64292 5540 64348
rect 5596 64292 8430 64348
rect 8486 64292 10740 64348
rect 5284 64288 10740 64292
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64348 16740 64352
rect 11284 64292 11320 64348
rect 11376 64292 14210 64348
rect 14266 64292 16740 64348
rect 11284 64288 16740 64292
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64348 17140 64352
rect 17124 64288 17140 64292
rect 17204 64288 17220 64352
rect 17284 64348 22740 64352
rect 17284 64292 19990 64348
rect 20046 64292 22740 64348
rect 17284 64288 22740 64292
rect 22804 64288 22820 64352
rect 22884 64348 22900 64352
rect 22884 64288 22900 64292
rect 22964 64288 22980 64352
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64348 28740 64352
rect 23284 64292 25770 64348
rect 25826 64292 28660 64348
rect 28716 64292 28740 64348
rect 23284 64288 28740 64292
rect 28804 64288 28820 64352
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64348 34740 64352
rect 29284 64292 31550 64348
rect 31606 64292 34440 64348
rect 34496 64292 34740 64348
rect 29284 64288 34740 64292
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64348 40740 64352
rect 35284 64292 37330 64348
rect 37386 64292 40220 64348
rect 40276 64292 40740 64348
rect 35284 64288 40740 64292
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64348 46740 64352
rect 41284 64292 43110 64348
rect 43166 64292 46000 64348
rect 46056 64292 46740 64348
rect 41284 64288 46740 64292
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64348 52740 64352
rect 47284 64292 49008 64348
rect 49064 64292 52237 64348
rect 52293 64292 52740 64348
rect 47284 64288 52740 64292
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64348 58740 64352
rect 53284 64292 53638 64348
rect 53694 64292 53806 64348
rect 53862 64292 54550 64348
rect 54606 64292 54940 64348
rect 54996 64292 55656 64348
rect 55712 64292 56234 64348
rect 56290 64292 56679 64348
rect 56735 64292 56983 64348
rect 57039 64292 57825 64348
rect 57881 64292 58465 64348
rect 58521 64292 58740 64348
rect 53284 64288 58740 64292
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64348 59060 64352
rect 59044 64292 59048 64348
rect 59044 64288 59060 64292
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64348 64740 64352
rect 59284 64292 60326 64348
rect 60382 64292 60484 64348
rect 60540 64292 62528 64348
rect 62584 64292 62608 64348
rect 62664 64292 64740 64348
rect 59284 64288 64740 64292
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64348 75028 64352
rect 71284 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 75028 64348
rect 71284 64288 75028 64292
rect 964 64264 75028 64288
rect 964 62240 75028 62264
rect 964 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62236 2220 62240
rect 2284 62236 7740 62240
rect 2320 62180 5393 62236
rect 5449 62180 7740 62236
rect 2204 62176 2220 62180
rect 2284 62176 7740 62180
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62236 13740 62240
rect 8339 62180 11173 62236
rect 11229 62180 13740 62236
rect 8284 62176 13740 62180
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62176 14220 62240
rect 14284 62236 19740 62240
rect 14284 62180 16953 62236
rect 17009 62180 19740 62236
rect 14284 62176 19740 62180
rect 19804 62176 19820 62240
rect 19884 62236 19900 62240
rect 19899 62180 19900 62236
rect 19884 62176 19900 62180
rect 19964 62176 19980 62240
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62236 25740 62240
rect 20284 62180 22733 62236
rect 22789 62180 25623 62236
rect 25679 62180 25740 62236
rect 20284 62176 25740 62180
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62236 31740 62240
rect 26284 62180 28513 62236
rect 28569 62180 31403 62236
rect 31459 62180 31740 62236
rect 26284 62176 31740 62180
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62236 37740 62240
rect 32284 62180 34293 62236
rect 34349 62180 37183 62236
rect 37239 62180 37740 62236
rect 32284 62176 37740 62180
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62236 43740 62240
rect 38284 62180 40073 62236
rect 40129 62180 42963 62236
rect 43019 62180 43740 62236
rect 38284 62176 43740 62180
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62236 49740 62240
rect 44284 62180 45853 62236
rect 45909 62180 48800 62236
rect 48856 62180 49662 62236
rect 49718 62180 49740 62236
rect 44284 62176 49740 62180
rect 49804 62176 49820 62240
rect 49884 62176 49900 62240
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62236 55740 62240
rect 50284 62180 52956 62236
rect 53012 62180 53114 62236
rect 53170 62180 53470 62236
rect 53526 62180 54788 62236
rect 54844 62180 55381 62236
rect 55437 62180 55740 62236
rect 50284 62176 55740 62180
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62236 61740 62240
rect 56284 62180 56527 62236
rect 56583 62180 57963 62236
rect 58019 62180 58043 62236
rect 58099 62180 59206 62236
rect 59262 62180 59364 62236
rect 59420 62180 59672 62236
rect 59728 62180 59818 62236
rect 59874 62180 59954 62236
rect 60010 62180 60034 62236
rect 60090 62180 61740 62236
rect 56284 62176 61740 62180
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62236 67740 62240
rect 62284 62180 62326 62236
rect 62382 62180 62406 62236
rect 62462 62180 67740 62236
rect 62284 62176 67740 62180
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62236 73740 62240
rect 68284 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 73740 62236
rect 68284 62176 73740 62180
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 75028 62240
rect 964 62160 75028 62176
rect 964 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62156 2220 62160
rect 2284 62156 7740 62160
rect 2320 62100 5393 62156
rect 5449 62100 7740 62156
rect 2204 62096 2220 62100
rect 2284 62096 7740 62100
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62156 13740 62160
rect 8339 62100 11173 62156
rect 11229 62100 13740 62156
rect 8284 62096 13740 62100
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62096 14220 62160
rect 14284 62156 19740 62160
rect 14284 62100 16953 62156
rect 17009 62100 19740 62156
rect 14284 62096 19740 62100
rect 19804 62096 19820 62160
rect 19884 62156 19900 62160
rect 19899 62100 19900 62156
rect 19884 62096 19900 62100
rect 19964 62096 19980 62160
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62156 25740 62160
rect 20284 62100 22733 62156
rect 22789 62100 25623 62156
rect 25679 62100 25740 62156
rect 20284 62096 25740 62100
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62156 31740 62160
rect 26284 62100 28513 62156
rect 28569 62100 31403 62156
rect 31459 62100 31740 62156
rect 26284 62096 31740 62100
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62156 37740 62160
rect 32284 62100 34293 62156
rect 34349 62100 37183 62156
rect 37239 62100 37740 62156
rect 32284 62096 37740 62100
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62156 43740 62160
rect 38284 62100 40073 62156
rect 40129 62100 42963 62156
rect 43019 62100 43740 62156
rect 38284 62096 43740 62100
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62156 49740 62160
rect 44284 62100 45853 62156
rect 45909 62100 48800 62156
rect 48856 62100 49662 62156
rect 49718 62100 49740 62156
rect 44284 62096 49740 62100
rect 49804 62096 49820 62160
rect 49884 62096 49900 62160
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62156 55740 62160
rect 50284 62100 52956 62156
rect 53012 62100 53114 62156
rect 53170 62100 53470 62156
rect 53526 62100 54788 62156
rect 54844 62100 55381 62156
rect 55437 62100 55740 62156
rect 50284 62096 55740 62100
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62156 61740 62160
rect 56284 62100 56527 62156
rect 56583 62100 57963 62156
rect 58019 62100 58043 62156
rect 58099 62100 59206 62156
rect 59262 62100 59364 62156
rect 59420 62100 59672 62156
rect 59728 62100 59818 62156
rect 59874 62100 59954 62156
rect 60010 62100 60034 62156
rect 60090 62100 61740 62156
rect 56284 62096 61740 62100
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62156 67740 62160
rect 62284 62100 62326 62156
rect 62382 62100 62406 62156
rect 62462 62100 67740 62156
rect 62284 62096 67740 62100
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62156 73740 62160
rect 68284 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 73740 62156
rect 68284 62096 73740 62100
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 75028 62160
rect 964 62080 75028 62096
rect 964 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62076 2220 62080
rect 2284 62076 7740 62080
rect 2320 62020 5393 62076
rect 5449 62020 7740 62076
rect 2204 62016 2220 62020
rect 2284 62016 7740 62020
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62076 13740 62080
rect 8339 62020 11173 62076
rect 11229 62020 13740 62076
rect 8284 62016 13740 62020
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62016 14220 62080
rect 14284 62076 19740 62080
rect 14284 62020 16953 62076
rect 17009 62020 19740 62076
rect 14284 62016 19740 62020
rect 19804 62016 19820 62080
rect 19884 62076 19900 62080
rect 19899 62020 19900 62076
rect 19884 62016 19900 62020
rect 19964 62016 19980 62080
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62076 25740 62080
rect 20284 62020 22733 62076
rect 22789 62020 25623 62076
rect 25679 62020 25740 62076
rect 20284 62016 25740 62020
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62076 31740 62080
rect 26284 62020 28513 62076
rect 28569 62020 31403 62076
rect 31459 62020 31740 62076
rect 26284 62016 31740 62020
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62076 37740 62080
rect 32284 62020 34293 62076
rect 34349 62020 37183 62076
rect 37239 62020 37740 62076
rect 32284 62016 37740 62020
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62076 43740 62080
rect 38284 62020 40073 62076
rect 40129 62020 42963 62076
rect 43019 62020 43740 62076
rect 38284 62016 43740 62020
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62076 49740 62080
rect 44284 62020 45853 62076
rect 45909 62020 48800 62076
rect 48856 62020 49662 62076
rect 49718 62020 49740 62076
rect 44284 62016 49740 62020
rect 49804 62016 49820 62080
rect 49884 62016 49900 62080
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62076 55740 62080
rect 50284 62020 52956 62076
rect 53012 62020 53114 62076
rect 53170 62020 53470 62076
rect 53526 62020 54788 62076
rect 54844 62020 55381 62076
rect 55437 62020 55740 62076
rect 50284 62016 55740 62020
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62076 61740 62080
rect 56284 62020 56527 62076
rect 56583 62020 57963 62076
rect 58019 62020 58043 62076
rect 58099 62020 59206 62076
rect 59262 62020 59364 62076
rect 59420 62020 59672 62076
rect 59728 62020 59818 62076
rect 59874 62020 59954 62076
rect 60010 62020 60034 62076
rect 60090 62020 61740 62076
rect 56284 62016 61740 62020
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62076 67740 62080
rect 62284 62020 62326 62076
rect 62382 62020 62406 62076
rect 62462 62020 67740 62076
rect 62284 62016 67740 62020
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62076 73740 62080
rect 68284 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 73740 62076
rect 68284 62016 73740 62020
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 75028 62080
rect 964 62000 75028 62016
rect 964 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61996 2220 62000
rect 2284 61996 7740 62000
rect 2320 61940 5393 61996
rect 5449 61940 7740 61996
rect 2204 61936 2220 61940
rect 2284 61936 7740 61940
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61996 13740 62000
rect 8339 61940 11173 61996
rect 11229 61940 13740 61996
rect 8284 61936 13740 61940
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61936 14220 62000
rect 14284 61996 19740 62000
rect 14284 61940 16953 61996
rect 17009 61940 19740 61996
rect 14284 61936 19740 61940
rect 19804 61936 19820 62000
rect 19884 61996 19900 62000
rect 19899 61940 19900 61996
rect 19884 61936 19900 61940
rect 19964 61936 19980 62000
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61996 25740 62000
rect 20284 61940 22733 61996
rect 22789 61940 25623 61996
rect 25679 61940 25740 61996
rect 20284 61936 25740 61940
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61996 31740 62000
rect 26284 61940 28513 61996
rect 28569 61940 31403 61996
rect 31459 61940 31740 61996
rect 26284 61936 31740 61940
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61996 37740 62000
rect 32284 61940 34293 61996
rect 34349 61940 37183 61996
rect 37239 61940 37740 61996
rect 32284 61936 37740 61940
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61996 43740 62000
rect 38284 61940 40073 61996
rect 40129 61940 42963 61996
rect 43019 61940 43740 61996
rect 38284 61936 43740 61940
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61996 49740 62000
rect 44284 61940 45853 61996
rect 45909 61940 48800 61996
rect 48856 61940 49662 61996
rect 49718 61940 49740 61996
rect 44284 61936 49740 61940
rect 49804 61936 49820 62000
rect 49884 61936 49900 62000
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61996 55740 62000
rect 50284 61940 52956 61996
rect 53012 61940 53114 61996
rect 53170 61940 53470 61996
rect 53526 61940 54788 61996
rect 54844 61940 55381 61996
rect 55437 61940 55740 61996
rect 50284 61936 55740 61940
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61996 61740 62000
rect 56284 61940 56527 61996
rect 56583 61940 57963 61996
rect 58019 61940 58043 61996
rect 58099 61940 59206 61996
rect 59262 61940 59364 61996
rect 59420 61940 59672 61996
rect 59728 61940 59818 61996
rect 59874 61940 59954 61996
rect 60010 61940 60034 61996
rect 60090 61940 61740 61996
rect 56284 61936 61740 61940
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61996 67740 62000
rect 62284 61940 62326 61996
rect 62382 61940 62406 61996
rect 62462 61940 67740 61996
rect 62284 61936 67740 61940
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61996 73740 62000
rect 68284 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 73740 61996
rect 68284 61936 73740 61940
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 75028 62000
rect 964 61912 75028 61936
rect 964 54592 75028 54616
rect 964 54588 4740 54592
rect 964 54532 2044 54588
rect 2100 54532 4740 54588
rect 964 54528 4740 54532
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54588 10740 54592
rect 5284 54532 5540 54588
rect 5596 54532 8430 54588
rect 8486 54532 10740 54588
rect 5284 54528 10740 54532
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54588 16740 54592
rect 11284 54532 11320 54588
rect 11376 54532 14210 54588
rect 14266 54532 16740 54588
rect 11284 54528 16740 54532
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54588 17140 54592
rect 17124 54528 17140 54532
rect 17204 54528 17220 54592
rect 17284 54588 22740 54592
rect 17284 54532 19990 54588
rect 20046 54532 22740 54588
rect 17284 54528 22740 54532
rect 22804 54528 22820 54592
rect 22884 54588 22900 54592
rect 22884 54528 22900 54532
rect 22964 54528 22980 54592
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54588 28740 54592
rect 23284 54532 25770 54588
rect 25826 54532 28660 54588
rect 28716 54532 28740 54588
rect 23284 54528 28740 54532
rect 28804 54528 28820 54592
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54588 34740 54592
rect 29284 54532 31550 54588
rect 31606 54532 34440 54588
rect 34496 54532 34740 54588
rect 29284 54528 34740 54532
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54588 40740 54592
rect 35284 54532 37330 54588
rect 37386 54532 40220 54588
rect 40276 54532 40740 54588
rect 35284 54528 40740 54532
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54588 46740 54592
rect 41284 54532 43110 54588
rect 43166 54532 46000 54588
rect 46056 54532 46740 54588
rect 41284 54528 46740 54532
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54588 52740 54592
rect 47284 54532 49008 54588
rect 49064 54532 52237 54588
rect 52293 54532 52740 54588
rect 47284 54528 52740 54532
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54588 58740 54592
rect 53284 54532 53638 54588
rect 53694 54532 53806 54588
rect 53862 54532 54550 54588
rect 54606 54532 54940 54588
rect 54996 54532 55656 54588
rect 55712 54532 56234 54588
rect 56290 54532 56679 54588
rect 56735 54532 56983 54588
rect 57039 54532 57825 54588
rect 57881 54532 58465 54588
rect 58521 54532 58740 54588
rect 53284 54528 58740 54532
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54588 59060 54592
rect 59044 54532 59048 54588
rect 59044 54528 59060 54532
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54588 64740 54592
rect 59284 54532 60326 54588
rect 60382 54532 60484 54588
rect 60540 54532 62528 54588
rect 62584 54532 62608 54588
rect 62664 54532 64740 54588
rect 59284 54528 64740 54532
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54588 75028 54592
rect 71284 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 75028 54588
rect 71284 54528 75028 54532
rect 964 54512 75028 54528
rect 964 54508 4740 54512
rect 964 54452 2044 54508
rect 2100 54452 4740 54508
rect 964 54448 4740 54452
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54508 10740 54512
rect 5284 54452 5540 54508
rect 5596 54452 8430 54508
rect 8486 54452 10740 54508
rect 5284 54448 10740 54452
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54508 16740 54512
rect 11284 54452 11320 54508
rect 11376 54452 14210 54508
rect 14266 54452 16740 54508
rect 11284 54448 16740 54452
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54508 17140 54512
rect 17124 54448 17140 54452
rect 17204 54448 17220 54512
rect 17284 54508 22740 54512
rect 17284 54452 19990 54508
rect 20046 54452 22740 54508
rect 17284 54448 22740 54452
rect 22804 54448 22820 54512
rect 22884 54508 22900 54512
rect 22884 54448 22900 54452
rect 22964 54448 22980 54512
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54508 28740 54512
rect 23284 54452 25770 54508
rect 25826 54452 28660 54508
rect 28716 54452 28740 54508
rect 23284 54448 28740 54452
rect 28804 54448 28820 54512
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54508 34740 54512
rect 29284 54452 31550 54508
rect 31606 54452 34440 54508
rect 34496 54452 34740 54508
rect 29284 54448 34740 54452
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54508 40740 54512
rect 35284 54452 37330 54508
rect 37386 54452 40220 54508
rect 40276 54452 40740 54508
rect 35284 54448 40740 54452
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54508 46740 54512
rect 41284 54452 43110 54508
rect 43166 54452 46000 54508
rect 46056 54452 46740 54508
rect 41284 54448 46740 54452
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54508 52740 54512
rect 47284 54452 49008 54508
rect 49064 54452 52237 54508
rect 52293 54452 52740 54508
rect 47284 54448 52740 54452
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54508 58740 54512
rect 53284 54452 53638 54508
rect 53694 54452 53806 54508
rect 53862 54452 54550 54508
rect 54606 54452 54940 54508
rect 54996 54452 55656 54508
rect 55712 54452 56234 54508
rect 56290 54452 56679 54508
rect 56735 54452 56983 54508
rect 57039 54452 57825 54508
rect 57881 54452 58465 54508
rect 58521 54452 58740 54508
rect 53284 54448 58740 54452
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54508 59060 54512
rect 59044 54452 59048 54508
rect 59044 54448 59060 54452
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54508 64740 54512
rect 59284 54452 60326 54508
rect 60382 54452 60484 54508
rect 60540 54452 62528 54508
rect 62584 54452 62608 54508
rect 62664 54452 64740 54508
rect 59284 54448 64740 54452
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54508 75028 54512
rect 71284 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 75028 54508
rect 71284 54448 75028 54452
rect 964 54432 75028 54448
rect 964 54428 4740 54432
rect 964 54372 2044 54428
rect 2100 54372 4740 54428
rect 964 54368 4740 54372
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54428 10740 54432
rect 5284 54372 5540 54428
rect 5596 54372 8430 54428
rect 8486 54372 10740 54428
rect 5284 54368 10740 54372
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54428 16740 54432
rect 11284 54372 11320 54428
rect 11376 54372 14210 54428
rect 14266 54372 16740 54428
rect 11284 54368 16740 54372
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54428 17140 54432
rect 17124 54368 17140 54372
rect 17204 54368 17220 54432
rect 17284 54428 22740 54432
rect 17284 54372 19990 54428
rect 20046 54372 22740 54428
rect 17284 54368 22740 54372
rect 22804 54368 22820 54432
rect 22884 54428 22900 54432
rect 22884 54368 22900 54372
rect 22964 54368 22980 54432
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54428 28740 54432
rect 23284 54372 25770 54428
rect 25826 54372 28660 54428
rect 28716 54372 28740 54428
rect 23284 54368 28740 54372
rect 28804 54368 28820 54432
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54428 34740 54432
rect 29284 54372 31550 54428
rect 31606 54372 34440 54428
rect 34496 54372 34740 54428
rect 29284 54368 34740 54372
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54428 40740 54432
rect 35284 54372 37330 54428
rect 37386 54372 40220 54428
rect 40276 54372 40740 54428
rect 35284 54368 40740 54372
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54428 46740 54432
rect 41284 54372 43110 54428
rect 43166 54372 46000 54428
rect 46056 54372 46740 54428
rect 41284 54368 46740 54372
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54428 52740 54432
rect 47284 54372 49008 54428
rect 49064 54372 52237 54428
rect 52293 54372 52740 54428
rect 47284 54368 52740 54372
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54428 58740 54432
rect 53284 54372 53638 54428
rect 53694 54372 53806 54428
rect 53862 54372 54550 54428
rect 54606 54372 54940 54428
rect 54996 54372 55656 54428
rect 55712 54372 56234 54428
rect 56290 54372 56679 54428
rect 56735 54372 56983 54428
rect 57039 54372 57825 54428
rect 57881 54372 58465 54428
rect 58521 54372 58740 54428
rect 53284 54368 58740 54372
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54428 59060 54432
rect 59044 54372 59048 54428
rect 59044 54368 59060 54372
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54428 64740 54432
rect 59284 54372 60326 54428
rect 60382 54372 60484 54428
rect 60540 54372 62528 54428
rect 62584 54372 62608 54428
rect 62664 54372 64740 54428
rect 59284 54368 64740 54372
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54428 75028 54432
rect 71284 54372 74216 54428
rect 74272 54372 74296 54428
rect 74352 54372 74376 54428
rect 74432 54372 74456 54428
rect 74512 54372 75028 54428
rect 71284 54368 75028 54372
rect 964 54352 75028 54368
rect 964 54348 4740 54352
rect 964 54292 2044 54348
rect 2100 54292 4740 54348
rect 964 54288 4740 54292
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54348 10740 54352
rect 5284 54292 5540 54348
rect 5596 54292 8430 54348
rect 8486 54292 10740 54348
rect 5284 54288 10740 54292
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54348 16740 54352
rect 11284 54292 11320 54348
rect 11376 54292 14210 54348
rect 14266 54292 16740 54348
rect 11284 54288 16740 54292
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54348 17140 54352
rect 17124 54288 17140 54292
rect 17204 54288 17220 54352
rect 17284 54348 22740 54352
rect 17284 54292 19990 54348
rect 20046 54292 22740 54348
rect 17284 54288 22740 54292
rect 22804 54288 22820 54352
rect 22884 54348 22900 54352
rect 22884 54288 22900 54292
rect 22964 54288 22980 54352
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54348 28740 54352
rect 23284 54292 25770 54348
rect 25826 54292 28660 54348
rect 28716 54292 28740 54348
rect 23284 54288 28740 54292
rect 28804 54288 28820 54352
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54348 34740 54352
rect 29284 54292 31550 54348
rect 31606 54292 34440 54348
rect 34496 54292 34740 54348
rect 29284 54288 34740 54292
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54348 40740 54352
rect 35284 54292 37330 54348
rect 37386 54292 40220 54348
rect 40276 54292 40740 54348
rect 35284 54288 40740 54292
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54348 46740 54352
rect 41284 54292 43110 54348
rect 43166 54292 46000 54348
rect 46056 54292 46740 54348
rect 41284 54288 46740 54292
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54348 52740 54352
rect 47284 54292 49008 54348
rect 49064 54292 52237 54348
rect 52293 54292 52740 54348
rect 47284 54288 52740 54292
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54348 58740 54352
rect 53284 54292 53638 54348
rect 53694 54292 53806 54348
rect 53862 54292 54550 54348
rect 54606 54292 54940 54348
rect 54996 54292 55656 54348
rect 55712 54292 56234 54348
rect 56290 54292 56679 54348
rect 56735 54292 56983 54348
rect 57039 54292 57825 54348
rect 57881 54292 58465 54348
rect 58521 54292 58740 54348
rect 53284 54288 58740 54292
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54348 59060 54352
rect 59044 54292 59048 54348
rect 59044 54288 59060 54292
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54348 64740 54352
rect 59284 54292 60326 54348
rect 60382 54292 60484 54348
rect 60540 54292 62528 54348
rect 62584 54292 62608 54348
rect 62664 54292 64740 54348
rect 59284 54288 64740 54292
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54348 75028 54352
rect 71284 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 75028 54348
rect 71284 54288 75028 54292
rect 964 54264 75028 54288
rect 63769 52594 63835 52597
rect 64086 52594 64092 52596
rect 63769 52592 64092 52594
rect 63769 52536 63774 52592
rect 63830 52536 64092 52592
rect 63769 52534 64092 52536
rect 63769 52531 63835 52534
rect 64086 52532 64092 52534
rect 64156 52532 64162 52596
rect 964 52240 75028 52264
rect 964 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52236 2220 52240
rect 2284 52236 7740 52240
rect 2320 52180 5393 52236
rect 5449 52180 7740 52236
rect 2204 52176 2220 52180
rect 2284 52176 7740 52180
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52236 13740 52240
rect 8339 52180 11173 52236
rect 11229 52180 13740 52236
rect 8284 52176 13740 52180
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52176 14220 52240
rect 14284 52236 19740 52240
rect 14284 52180 16953 52236
rect 17009 52180 19740 52236
rect 14284 52176 19740 52180
rect 19804 52176 19820 52240
rect 19884 52236 19900 52240
rect 19899 52180 19900 52236
rect 19884 52176 19900 52180
rect 19964 52176 19980 52240
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52236 25740 52240
rect 20284 52180 22733 52236
rect 22789 52180 25623 52236
rect 25679 52180 25740 52236
rect 20284 52176 25740 52180
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52236 31740 52240
rect 26284 52180 28513 52236
rect 28569 52180 31403 52236
rect 31459 52180 31740 52236
rect 26284 52176 31740 52180
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52236 37740 52240
rect 32284 52180 34293 52236
rect 34349 52180 37183 52236
rect 37239 52180 37740 52236
rect 32284 52176 37740 52180
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52236 43740 52240
rect 38284 52180 40073 52236
rect 40129 52180 42963 52236
rect 43019 52180 43740 52236
rect 38284 52176 43740 52180
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52236 49740 52240
rect 44284 52180 45853 52236
rect 45909 52180 48800 52236
rect 48856 52180 49662 52236
rect 49718 52180 49740 52236
rect 44284 52176 49740 52180
rect 49804 52176 49820 52240
rect 49884 52176 49900 52240
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52236 55740 52240
rect 50284 52180 52956 52236
rect 53012 52180 53114 52236
rect 53170 52180 53470 52236
rect 53526 52180 54788 52236
rect 54844 52180 55381 52236
rect 55437 52180 55740 52236
rect 50284 52176 55740 52180
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52236 61740 52240
rect 56284 52180 56527 52236
rect 56583 52180 57963 52236
rect 58019 52180 58043 52236
rect 58099 52180 59206 52236
rect 59262 52180 59364 52236
rect 59420 52180 59672 52236
rect 59728 52180 59818 52236
rect 59874 52180 59954 52236
rect 60010 52180 60034 52236
rect 60090 52180 61740 52236
rect 56284 52176 61740 52180
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52236 67740 52240
rect 62284 52180 62326 52236
rect 62382 52180 62406 52236
rect 62462 52180 67740 52236
rect 62284 52176 67740 52180
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52236 73740 52240
rect 68284 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 73740 52236
rect 68284 52176 73740 52180
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 75028 52240
rect 964 52160 75028 52176
rect 964 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52156 2220 52160
rect 2284 52156 7740 52160
rect 2320 52100 5393 52156
rect 5449 52100 7740 52156
rect 2204 52096 2220 52100
rect 2284 52096 7740 52100
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52156 13740 52160
rect 8339 52100 11173 52156
rect 11229 52100 13740 52156
rect 8284 52096 13740 52100
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52096 14220 52160
rect 14284 52156 19740 52160
rect 14284 52100 16953 52156
rect 17009 52100 19740 52156
rect 14284 52096 19740 52100
rect 19804 52096 19820 52160
rect 19884 52156 19900 52160
rect 19899 52100 19900 52156
rect 19884 52096 19900 52100
rect 19964 52096 19980 52160
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52156 25740 52160
rect 20284 52100 22733 52156
rect 22789 52100 25623 52156
rect 25679 52100 25740 52156
rect 20284 52096 25740 52100
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52156 31740 52160
rect 26284 52100 28513 52156
rect 28569 52100 31403 52156
rect 31459 52100 31740 52156
rect 26284 52096 31740 52100
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52156 37740 52160
rect 32284 52100 34293 52156
rect 34349 52100 37183 52156
rect 37239 52100 37740 52156
rect 32284 52096 37740 52100
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52156 43740 52160
rect 38284 52100 40073 52156
rect 40129 52100 42963 52156
rect 43019 52100 43740 52156
rect 38284 52096 43740 52100
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52156 49740 52160
rect 44284 52100 45853 52156
rect 45909 52100 48800 52156
rect 48856 52100 49662 52156
rect 49718 52100 49740 52156
rect 44284 52096 49740 52100
rect 49804 52096 49820 52160
rect 49884 52096 49900 52160
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52156 55740 52160
rect 50284 52100 52956 52156
rect 53012 52100 53114 52156
rect 53170 52100 53470 52156
rect 53526 52100 54788 52156
rect 54844 52100 55381 52156
rect 55437 52100 55740 52156
rect 50284 52096 55740 52100
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52156 61740 52160
rect 56284 52100 56527 52156
rect 56583 52100 57963 52156
rect 58019 52100 58043 52156
rect 58099 52100 59206 52156
rect 59262 52100 59364 52156
rect 59420 52100 59672 52156
rect 59728 52100 59818 52156
rect 59874 52100 59954 52156
rect 60010 52100 60034 52156
rect 60090 52100 61740 52156
rect 56284 52096 61740 52100
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52156 67740 52160
rect 62284 52100 62326 52156
rect 62382 52100 62406 52156
rect 62462 52100 67740 52156
rect 62284 52096 67740 52100
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52156 73740 52160
rect 68284 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 73740 52156
rect 68284 52096 73740 52100
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 75028 52160
rect 964 52080 75028 52096
rect 964 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52076 2220 52080
rect 2284 52076 7740 52080
rect 2320 52020 5393 52076
rect 5449 52020 7740 52076
rect 2204 52016 2220 52020
rect 2284 52016 7740 52020
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52076 13740 52080
rect 8339 52020 11173 52076
rect 11229 52020 13740 52076
rect 8284 52016 13740 52020
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52016 14220 52080
rect 14284 52076 19740 52080
rect 14284 52020 16953 52076
rect 17009 52020 19740 52076
rect 14284 52016 19740 52020
rect 19804 52016 19820 52080
rect 19884 52076 19900 52080
rect 19899 52020 19900 52076
rect 19884 52016 19900 52020
rect 19964 52016 19980 52080
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52076 25740 52080
rect 20284 52020 22733 52076
rect 22789 52020 25623 52076
rect 25679 52020 25740 52076
rect 20284 52016 25740 52020
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52076 31740 52080
rect 26284 52020 28513 52076
rect 28569 52020 31403 52076
rect 31459 52020 31740 52076
rect 26284 52016 31740 52020
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52076 37740 52080
rect 32284 52020 34293 52076
rect 34349 52020 37183 52076
rect 37239 52020 37740 52076
rect 32284 52016 37740 52020
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52076 43740 52080
rect 38284 52020 40073 52076
rect 40129 52020 42963 52076
rect 43019 52020 43740 52076
rect 38284 52016 43740 52020
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52076 49740 52080
rect 44284 52020 45853 52076
rect 45909 52020 48800 52076
rect 48856 52020 49662 52076
rect 49718 52020 49740 52076
rect 44284 52016 49740 52020
rect 49804 52016 49820 52080
rect 49884 52016 49900 52080
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52076 55740 52080
rect 50284 52020 52956 52076
rect 53012 52020 53114 52076
rect 53170 52020 53470 52076
rect 53526 52020 54788 52076
rect 54844 52020 55381 52076
rect 55437 52020 55740 52076
rect 50284 52016 55740 52020
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52076 61740 52080
rect 56284 52020 56527 52076
rect 56583 52020 57963 52076
rect 58019 52020 58043 52076
rect 58099 52020 59206 52076
rect 59262 52020 59364 52076
rect 59420 52020 59672 52076
rect 59728 52020 59818 52076
rect 59874 52020 59954 52076
rect 60010 52020 60034 52076
rect 60090 52020 61740 52076
rect 56284 52016 61740 52020
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52076 67740 52080
rect 62284 52020 62326 52076
rect 62382 52020 62406 52076
rect 62462 52020 67740 52076
rect 62284 52016 67740 52020
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52076 73740 52080
rect 68284 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 73740 52076
rect 68284 52016 73740 52020
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 75028 52080
rect 964 52000 75028 52016
rect 964 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51996 2220 52000
rect 2284 51996 7740 52000
rect 2320 51940 5393 51996
rect 5449 51940 7740 51996
rect 2204 51936 2220 51940
rect 2284 51936 7740 51940
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51996 13740 52000
rect 8339 51940 11173 51996
rect 11229 51940 13740 51996
rect 8284 51936 13740 51940
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51936 14220 52000
rect 14284 51996 19740 52000
rect 14284 51940 16953 51996
rect 17009 51940 19740 51996
rect 14284 51936 19740 51940
rect 19804 51936 19820 52000
rect 19884 51996 19900 52000
rect 19899 51940 19900 51996
rect 19884 51936 19900 51940
rect 19964 51936 19980 52000
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51996 25740 52000
rect 20284 51940 22733 51996
rect 22789 51940 25623 51996
rect 25679 51940 25740 51996
rect 20284 51936 25740 51940
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51996 31740 52000
rect 26284 51940 28513 51996
rect 28569 51940 31403 51996
rect 31459 51940 31740 51996
rect 26284 51936 31740 51940
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51996 37740 52000
rect 32284 51940 34293 51996
rect 34349 51940 37183 51996
rect 37239 51940 37740 51996
rect 32284 51936 37740 51940
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51996 43740 52000
rect 38284 51940 40073 51996
rect 40129 51940 42963 51996
rect 43019 51940 43740 51996
rect 38284 51936 43740 51940
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51996 49740 52000
rect 44284 51940 45853 51996
rect 45909 51940 48800 51996
rect 48856 51940 49662 51996
rect 49718 51940 49740 51996
rect 44284 51936 49740 51940
rect 49804 51936 49820 52000
rect 49884 51936 49900 52000
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51996 55740 52000
rect 50284 51940 52956 51996
rect 53012 51940 53114 51996
rect 53170 51940 53470 51996
rect 53526 51940 54788 51996
rect 54844 51940 55381 51996
rect 55437 51940 55740 51996
rect 50284 51936 55740 51940
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51996 61740 52000
rect 56284 51940 56527 51996
rect 56583 51940 57963 51996
rect 58019 51940 58043 51996
rect 58099 51940 59206 51996
rect 59262 51940 59364 51996
rect 59420 51940 59672 51996
rect 59728 51940 59818 51996
rect 59874 51940 59954 51996
rect 60010 51940 60034 51996
rect 60090 51940 61740 51996
rect 56284 51936 61740 51940
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51996 67740 52000
rect 62284 51940 62326 51996
rect 62382 51940 62406 51996
rect 62462 51940 67740 51996
rect 62284 51936 67740 51940
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51996 73740 52000
rect 68284 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 73740 51996
rect 68284 51936 73740 51940
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 75028 52000
rect 964 51912 75028 51936
rect 63769 50282 63835 50285
rect 64270 50282 64276 50284
rect 63769 50280 64276 50282
rect 63769 50224 63774 50280
rect 63830 50224 64276 50280
rect 63769 50222 64276 50224
rect 63769 50219 63835 50222
rect 64270 50220 64276 50222
rect 64340 50220 64346 50284
rect 64965 48106 65031 48109
rect 65558 48106 65564 48108
rect 64965 48104 65564 48106
rect 64965 48048 64970 48104
rect 65026 48048 65564 48104
rect 64965 48046 65564 48048
rect 64965 48043 65031 48046
rect 65558 48044 65564 48046
rect 65628 48044 65634 48108
rect 64413 47700 64479 47701
rect 64413 47696 64460 47700
rect 64524 47698 64530 47700
rect 64413 47640 64418 47696
rect 64413 47636 64460 47640
rect 64524 47638 64570 47698
rect 64524 47636 64530 47638
rect 64413 47635 64479 47636
rect 63166 44780 63172 44844
rect 63236 44842 63242 44844
rect 65241 44842 65307 44845
rect 63236 44840 65307 44842
rect 63236 44784 65246 44840
rect 65302 44784 65307 44840
rect 63236 44782 65307 44784
rect 63236 44780 63242 44782
rect 65241 44779 65307 44782
rect 964 44592 75028 44616
rect 964 44588 4740 44592
rect 964 44532 2044 44588
rect 2100 44532 4740 44588
rect 964 44528 4740 44532
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44588 10740 44592
rect 5284 44532 5540 44588
rect 5596 44532 8430 44588
rect 8486 44532 10740 44588
rect 5284 44528 10740 44532
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44588 16740 44592
rect 11284 44532 11320 44588
rect 11376 44532 14210 44588
rect 14266 44532 16740 44588
rect 11284 44528 16740 44532
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44588 17140 44592
rect 17124 44528 17140 44532
rect 17204 44528 17220 44592
rect 17284 44588 22740 44592
rect 17284 44532 19990 44588
rect 20046 44532 22740 44588
rect 17284 44528 22740 44532
rect 22804 44528 22820 44592
rect 22884 44588 22900 44592
rect 22884 44528 22900 44532
rect 22964 44528 22980 44592
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44588 28740 44592
rect 23284 44532 25770 44588
rect 25826 44532 28660 44588
rect 28716 44532 28740 44588
rect 23284 44528 28740 44532
rect 28804 44528 28820 44592
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44588 34740 44592
rect 29284 44532 31550 44588
rect 31606 44532 34440 44588
rect 34496 44532 34740 44588
rect 29284 44528 34740 44532
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44588 40740 44592
rect 35284 44532 37330 44588
rect 37386 44532 40220 44588
rect 40276 44532 40740 44588
rect 35284 44528 40740 44532
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44588 46740 44592
rect 41284 44532 43110 44588
rect 43166 44532 46000 44588
rect 46056 44532 46740 44588
rect 41284 44528 46740 44532
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44588 52740 44592
rect 47284 44532 52237 44588
rect 52293 44532 52740 44588
rect 47284 44528 52740 44532
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44588 58740 44592
rect 53284 44532 53638 44588
rect 53694 44532 54550 44588
rect 54606 44532 54940 44588
rect 54996 44532 55656 44588
rect 55712 44532 56234 44588
rect 56290 44532 56679 44588
rect 56735 44532 56983 44588
rect 57039 44532 57825 44588
rect 57881 44532 58349 44588
rect 58405 44532 58740 44588
rect 53284 44528 58740 44532
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44588 59060 44592
rect 59044 44532 59048 44588
rect 59044 44528 59060 44532
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44588 64740 44592
rect 59284 44532 60326 44588
rect 60382 44532 60484 44588
rect 60540 44532 62528 44588
rect 62584 44532 62608 44588
rect 62664 44532 64740 44588
rect 59284 44528 64740 44532
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44588 75028 44592
rect 71284 44532 74216 44588
rect 74272 44532 74296 44588
rect 74352 44532 74376 44588
rect 74432 44532 74456 44588
rect 74512 44532 75028 44588
rect 71284 44528 75028 44532
rect 964 44512 75028 44528
rect 964 44508 4740 44512
rect 964 44452 2044 44508
rect 2100 44452 4740 44508
rect 964 44448 4740 44452
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44508 10740 44512
rect 5284 44452 5540 44508
rect 5596 44452 8430 44508
rect 8486 44452 10740 44508
rect 5284 44448 10740 44452
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44508 16740 44512
rect 11284 44452 11320 44508
rect 11376 44452 14210 44508
rect 14266 44452 16740 44508
rect 11284 44448 16740 44452
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44508 17140 44512
rect 17124 44448 17140 44452
rect 17204 44448 17220 44512
rect 17284 44508 22740 44512
rect 17284 44452 19990 44508
rect 20046 44452 22740 44508
rect 17284 44448 22740 44452
rect 22804 44448 22820 44512
rect 22884 44508 22900 44512
rect 22884 44448 22900 44452
rect 22964 44448 22980 44512
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44508 28740 44512
rect 23284 44452 25770 44508
rect 25826 44452 28660 44508
rect 28716 44452 28740 44508
rect 23284 44448 28740 44452
rect 28804 44448 28820 44512
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44508 34740 44512
rect 29284 44452 31550 44508
rect 31606 44452 34440 44508
rect 34496 44452 34740 44508
rect 29284 44448 34740 44452
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44508 40740 44512
rect 35284 44452 37330 44508
rect 37386 44452 40220 44508
rect 40276 44452 40740 44508
rect 35284 44448 40740 44452
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44508 46740 44512
rect 41284 44452 43110 44508
rect 43166 44452 46000 44508
rect 46056 44452 46740 44508
rect 41284 44448 46740 44452
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44508 52740 44512
rect 47284 44452 52237 44508
rect 52293 44452 52740 44508
rect 47284 44448 52740 44452
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44508 58740 44512
rect 53284 44452 53638 44508
rect 53694 44452 54550 44508
rect 54606 44452 54940 44508
rect 54996 44452 55656 44508
rect 55712 44452 56234 44508
rect 56290 44452 56679 44508
rect 56735 44452 56983 44508
rect 57039 44452 57825 44508
rect 57881 44452 58349 44508
rect 58405 44452 58740 44508
rect 53284 44448 58740 44452
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44508 59060 44512
rect 59044 44452 59048 44508
rect 59044 44448 59060 44452
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44508 64740 44512
rect 59284 44452 60326 44508
rect 60382 44452 60484 44508
rect 60540 44452 62528 44508
rect 62584 44452 62608 44508
rect 62664 44452 64740 44508
rect 59284 44448 64740 44452
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44508 75028 44512
rect 71284 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 75028 44508
rect 71284 44448 75028 44452
rect 964 44432 75028 44448
rect 964 44428 4740 44432
rect 964 44372 2044 44428
rect 2100 44372 4740 44428
rect 964 44368 4740 44372
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44428 10740 44432
rect 5284 44372 5540 44428
rect 5596 44372 8430 44428
rect 8486 44372 10740 44428
rect 5284 44368 10740 44372
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44428 16740 44432
rect 11284 44372 11320 44428
rect 11376 44372 14210 44428
rect 14266 44372 16740 44428
rect 11284 44368 16740 44372
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44428 17140 44432
rect 17124 44368 17140 44372
rect 17204 44368 17220 44432
rect 17284 44428 22740 44432
rect 17284 44372 19990 44428
rect 20046 44372 22740 44428
rect 17284 44368 22740 44372
rect 22804 44368 22820 44432
rect 22884 44428 22900 44432
rect 22884 44368 22900 44372
rect 22964 44368 22980 44432
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44428 28740 44432
rect 23284 44372 25770 44428
rect 25826 44372 28660 44428
rect 28716 44372 28740 44428
rect 23284 44368 28740 44372
rect 28804 44368 28820 44432
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44428 34740 44432
rect 29284 44372 31550 44428
rect 31606 44372 34440 44428
rect 34496 44372 34740 44428
rect 29284 44368 34740 44372
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44428 40740 44432
rect 35284 44372 37330 44428
rect 37386 44372 40220 44428
rect 40276 44372 40740 44428
rect 35284 44368 40740 44372
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44428 46740 44432
rect 41284 44372 43110 44428
rect 43166 44372 46000 44428
rect 46056 44372 46740 44428
rect 41284 44368 46740 44372
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44428 52740 44432
rect 47284 44372 52237 44428
rect 52293 44372 52740 44428
rect 47284 44368 52740 44372
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44428 58740 44432
rect 53284 44372 53638 44428
rect 53694 44372 54550 44428
rect 54606 44372 54940 44428
rect 54996 44372 55656 44428
rect 55712 44372 56234 44428
rect 56290 44372 56679 44428
rect 56735 44372 56983 44428
rect 57039 44372 57825 44428
rect 57881 44372 58349 44428
rect 58405 44372 58740 44428
rect 53284 44368 58740 44372
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44428 59060 44432
rect 59044 44372 59048 44428
rect 59044 44368 59060 44372
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44428 64740 44432
rect 59284 44372 60326 44428
rect 60382 44372 60484 44428
rect 60540 44372 62528 44428
rect 62584 44372 62608 44428
rect 62664 44372 64740 44428
rect 59284 44368 64740 44372
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44428 75028 44432
rect 71284 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 75028 44428
rect 71284 44368 75028 44372
rect 964 44352 75028 44368
rect 964 44348 4740 44352
rect 964 44292 2044 44348
rect 2100 44292 4740 44348
rect 964 44288 4740 44292
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44348 10740 44352
rect 5284 44292 5540 44348
rect 5596 44292 8430 44348
rect 8486 44292 10740 44348
rect 5284 44288 10740 44292
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44348 16740 44352
rect 11284 44292 11320 44348
rect 11376 44292 14210 44348
rect 14266 44292 16740 44348
rect 11284 44288 16740 44292
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44348 17140 44352
rect 17124 44288 17140 44292
rect 17204 44288 17220 44352
rect 17284 44348 22740 44352
rect 17284 44292 19990 44348
rect 20046 44292 22740 44348
rect 17284 44288 22740 44292
rect 22804 44288 22820 44352
rect 22884 44348 22900 44352
rect 22884 44288 22900 44292
rect 22964 44288 22980 44352
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44348 28740 44352
rect 23284 44292 25770 44348
rect 25826 44292 28660 44348
rect 28716 44292 28740 44348
rect 23284 44288 28740 44292
rect 28804 44288 28820 44352
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44348 34740 44352
rect 29284 44292 31550 44348
rect 31606 44292 34440 44348
rect 34496 44292 34740 44348
rect 29284 44288 34740 44292
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44348 40740 44352
rect 35284 44292 37330 44348
rect 37386 44292 40220 44348
rect 40276 44292 40740 44348
rect 35284 44288 40740 44292
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44348 46740 44352
rect 41284 44292 43110 44348
rect 43166 44292 46000 44348
rect 46056 44292 46740 44348
rect 41284 44288 46740 44292
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44348 52740 44352
rect 47284 44292 52237 44348
rect 52293 44292 52740 44348
rect 47284 44288 52740 44292
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44348 58740 44352
rect 53284 44292 53638 44348
rect 53694 44292 54550 44348
rect 54606 44292 54940 44348
rect 54996 44292 55656 44348
rect 55712 44292 56234 44348
rect 56290 44292 56679 44348
rect 56735 44292 56983 44348
rect 57039 44292 57825 44348
rect 57881 44292 58349 44348
rect 58405 44292 58740 44348
rect 53284 44288 58740 44292
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44348 59060 44352
rect 59044 44292 59048 44348
rect 59044 44288 59060 44292
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44348 64740 44352
rect 59284 44292 60326 44348
rect 60382 44292 60484 44348
rect 60540 44292 62528 44348
rect 62584 44292 62608 44348
rect 62664 44292 64740 44348
rect 59284 44288 64740 44292
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44348 75028 44352
rect 71284 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 75028 44348
rect 71284 44288 75028 44292
rect 964 44264 75028 44288
rect 63769 43346 63835 43349
rect 63902 43346 63908 43348
rect 63769 43344 63908 43346
rect 63769 43288 63774 43344
rect 63830 43288 63908 43344
rect 63769 43286 63908 43288
rect 63769 43283 63835 43286
rect 63902 43284 63908 43286
rect 63972 43284 63978 43348
rect 964 42240 75028 42264
rect 964 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42236 2220 42240
rect 2284 42236 7740 42240
rect 2320 42180 5393 42236
rect 5449 42180 7740 42236
rect 2204 42176 2220 42180
rect 2284 42176 7740 42180
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42236 13740 42240
rect 8339 42180 11173 42236
rect 11229 42180 13740 42236
rect 8284 42176 13740 42180
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42176 14220 42240
rect 14284 42236 19740 42240
rect 14284 42180 16953 42236
rect 17009 42180 19740 42236
rect 14284 42176 19740 42180
rect 19804 42176 19820 42240
rect 19884 42236 19900 42240
rect 19899 42180 19900 42236
rect 19884 42176 19900 42180
rect 19964 42176 19980 42240
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42236 25740 42240
rect 20284 42180 22733 42236
rect 22789 42180 25623 42236
rect 25679 42180 25740 42236
rect 20284 42176 25740 42180
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42236 31740 42240
rect 26284 42180 28513 42236
rect 28569 42180 31403 42236
rect 31459 42180 31740 42236
rect 26284 42176 31740 42180
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42236 37740 42240
rect 32284 42180 34293 42236
rect 34349 42180 37183 42236
rect 37239 42180 37740 42236
rect 32284 42176 37740 42180
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42236 43740 42240
rect 38284 42180 40073 42236
rect 40129 42180 42963 42236
rect 43019 42180 43740 42236
rect 38284 42176 43740 42180
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42236 49740 42240
rect 44284 42180 45853 42236
rect 45909 42180 48800 42236
rect 48856 42180 49662 42236
rect 49718 42180 49740 42236
rect 44284 42176 49740 42180
rect 49804 42176 49820 42240
rect 49884 42176 49900 42240
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42236 55740 42240
rect 50284 42180 52956 42236
rect 53012 42180 53114 42236
rect 53170 42180 53470 42236
rect 53526 42180 54788 42236
rect 54844 42180 55381 42236
rect 55437 42180 55740 42236
rect 50284 42176 55740 42180
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42236 61740 42240
rect 56284 42180 56527 42236
rect 56583 42180 57963 42236
rect 58019 42180 58043 42236
rect 58099 42180 59206 42236
rect 59262 42180 59364 42236
rect 59420 42180 59672 42236
rect 59728 42180 59818 42236
rect 59874 42180 59954 42236
rect 60010 42180 60034 42236
rect 60090 42180 61740 42236
rect 56284 42176 61740 42180
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42236 67740 42240
rect 62284 42180 62326 42236
rect 62382 42180 62406 42236
rect 62462 42180 67740 42236
rect 62284 42176 67740 42180
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42236 73740 42240
rect 68284 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 73740 42236
rect 68284 42176 73740 42180
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 75028 42240
rect 964 42160 75028 42176
rect 964 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42156 2220 42160
rect 2284 42156 7740 42160
rect 2320 42100 5393 42156
rect 5449 42100 7740 42156
rect 2204 42096 2220 42100
rect 2284 42096 7740 42100
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42156 13740 42160
rect 8339 42100 11173 42156
rect 11229 42100 13740 42156
rect 8284 42096 13740 42100
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42096 14220 42160
rect 14284 42156 19740 42160
rect 14284 42100 16953 42156
rect 17009 42100 19740 42156
rect 14284 42096 19740 42100
rect 19804 42096 19820 42160
rect 19884 42156 19900 42160
rect 19899 42100 19900 42156
rect 19884 42096 19900 42100
rect 19964 42096 19980 42160
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42156 25740 42160
rect 20284 42100 22733 42156
rect 22789 42100 25623 42156
rect 25679 42100 25740 42156
rect 20284 42096 25740 42100
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42156 31740 42160
rect 26284 42100 28513 42156
rect 28569 42100 31403 42156
rect 31459 42100 31740 42156
rect 26284 42096 31740 42100
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42156 37740 42160
rect 32284 42100 34293 42156
rect 34349 42100 37183 42156
rect 37239 42100 37740 42156
rect 32284 42096 37740 42100
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42156 43740 42160
rect 38284 42100 40073 42156
rect 40129 42100 42963 42156
rect 43019 42100 43740 42156
rect 38284 42096 43740 42100
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42156 49740 42160
rect 44284 42100 45853 42156
rect 45909 42100 48800 42156
rect 48856 42100 49662 42156
rect 49718 42100 49740 42156
rect 44284 42096 49740 42100
rect 49804 42096 49820 42160
rect 49884 42096 49900 42160
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42156 55740 42160
rect 50284 42100 52956 42156
rect 53012 42100 53114 42156
rect 53170 42100 53470 42156
rect 53526 42100 54788 42156
rect 54844 42100 55381 42156
rect 55437 42100 55740 42156
rect 50284 42096 55740 42100
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42156 61740 42160
rect 56284 42100 56527 42156
rect 56583 42100 57963 42156
rect 58019 42100 58043 42156
rect 58099 42100 59206 42156
rect 59262 42100 59364 42156
rect 59420 42100 59672 42156
rect 59728 42100 59818 42156
rect 59874 42100 59954 42156
rect 60010 42100 60034 42156
rect 60090 42100 61740 42156
rect 56284 42096 61740 42100
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42156 67740 42160
rect 62284 42100 62326 42156
rect 62382 42100 62406 42156
rect 62462 42100 67740 42156
rect 62284 42096 67740 42100
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42156 73740 42160
rect 68284 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 73740 42156
rect 68284 42096 73740 42100
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 75028 42160
rect 964 42080 75028 42096
rect 964 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42076 2220 42080
rect 2284 42076 7740 42080
rect 2320 42020 5393 42076
rect 5449 42020 7740 42076
rect 2204 42016 2220 42020
rect 2284 42016 7740 42020
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42076 13740 42080
rect 8339 42020 11173 42076
rect 11229 42020 13740 42076
rect 8284 42016 13740 42020
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42016 14220 42080
rect 14284 42076 19740 42080
rect 14284 42020 16953 42076
rect 17009 42020 19740 42076
rect 14284 42016 19740 42020
rect 19804 42016 19820 42080
rect 19884 42076 19900 42080
rect 19899 42020 19900 42076
rect 19884 42016 19900 42020
rect 19964 42016 19980 42080
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42076 25740 42080
rect 20284 42020 22733 42076
rect 22789 42020 25623 42076
rect 25679 42020 25740 42076
rect 20284 42016 25740 42020
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42076 31740 42080
rect 26284 42020 28513 42076
rect 28569 42020 31403 42076
rect 31459 42020 31740 42076
rect 26284 42016 31740 42020
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42076 37740 42080
rect 32284 42020 34293 42076
rect 34349 42020 37183 42076
rect 37239 42020 37740 42076
rect 32284 42016 37740 42020
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42076 43740 42080
rect 38284 42020 40073 42076
rect 40129 42020 42963 42076
rect 43019 42020 43740 42076
rect 38284 42016 43740 42020
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42076 49740 42080
rect 44284 42020 45853 42076
rect 45909 42020 48800 42076
rect 48856 42020 49662 42076
rect 49718 42020 49740 42076
rect 44284 42016 49740 42020
rect 49804 42016 49820 42080
rect 49884 42016 49900 42080
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42076 55740 42080
rect 50284 42020 52956 42076
rect 53012 42020 53114 42076
rect 53170 42020 53470 42076
rect 53526 42020 54788 42076
rect 54844 42020 55381 42076
rect 55437 42020 55740 42076
rect 50284 42016 55740 42020
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42076 61740 42080
rect 56284 42020 56527 42076
rect 56583 42020 57963 42076
rect 58019 42020 58043 42076
rect 58099 42020 59206 42076
rect 59262 42020 59364 42076
rect 59420 42020 59672 42076
rect 59728 42020 59818 42076
rect 59874 42020 59954 42076
rect 60010 42020 60034 42076
rect 60090 42020 61740 42076
rect 56284 42016 61740 42020
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42076 67740 42080
rect 62284 42020 62326 42076
rect 62382 42020 62406 42076
rect 62462 42020 67740 42076
rect 62284 42016 67740 42020
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42076 73740 42080
rect 68284 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 73740 42076
rect 68284 42016 73740 42020
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 75028 42080
rect 964 42000 75028 42016
rect 964 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41996 2220 42000
rect 2284 41996 7740 42000
rect 2320 41940 5393 41996
rect 5449 41940 7740 41996
rect 2204 41936 2220 41940
rect 2284 41936 7740 41940
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41996 13740 42000
rect 8339 41940 11173 41996
rect 11229 41940 13740 41996
rect 8284 41936 13740 41940
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41936 14220 42000
rect 14284 41996 19740 42000
rect 14284 41940 16953 41996
rect 17009 41940 19740 41996
rect 14284 41936 19740 41940
rect 19804 41936 19820 42000
rect 19884 41996 19900 42000
rect 19899 41940 19900 41996
rect 19884 41936 19900 41940
rect 19964 41936 19980 42000
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41996 25740 42000
rect 20284 41940 22733 41996
rect 22789 41940 25623 41996
rect 25679 41940 25740 41996
rect 20284 41936 25740 41940
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41996 31740 42000
rect 26284 41940 28513 41996
rect 28569 41940 31403 41996
rect 31459 41940 31740 41996
rect 26284 41936 31740 41940
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41996 37740 42000
rect 32284 41940 34293 41996
rect 34349 41940 37183 41996
rect 37239 41940 37740 41996
rect 32284 41936 37740 41940
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41996 43740 42000
rect 38284 41940 40073 41996
rect 40129 41940 42963 41996
rect 43019 41940 43740 41996
rect 38284 41936 43740 41940
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41996 49740 42000
rect 44284 41940 45853 41996
rect 45909 41940 48800 41996
rect 48856 41940 49662 41996
rect 49718 41940 49740 41996
rect 44284 41936 49740 41940
rect 49804 41936 49820 42000
rect 49884 41936 49900 42000
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41996 55740 42000
rect 50284 41940 52956 41996
rect 53012 41940 53114 41996
rect 53170 41940 53470 41996
rect 53526 41940 54788 41996
rect 54844 41940 55381 41996
rect 55437 41940 55740 41996
rect 50284 41936 55740 41940
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41996 61740 42000
rect 56284 41940 56527 41996
rect 56583 41940 57963 41996
rect 58019 41940 58043 41996
rect 58099 41940 59206 41996
rect 59262 41940 59364 41996
rect 59420 41940 59672 41996
rect 59728 41940 59818 41996
rect 59874 41940 59954 41996
rect 60010 41940 60034 41996
rect 60090 41940 61740 41996
rect 56284 41936 61740 41940
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41996 67740 42000
rect 62284 41940 62326 41996
rect 62382 41940 62406 41996
rect 62462 41940 67740 41996
rect 62284 41936 67740 41940
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41996 73740 42000
rect 68284 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 73740 41996
rect 68284 41936 73740 41940
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 75028 42000
rect 964 41912 75028 41936
rect 65241 40898 65307 40901
rect 65742 40898 65748 40900
rect 65241 40896 65748 40898
rect 65241 40840 65246 40896
rect 65302 40840 65748 40896
rect 65241 40838 65748 40840
rect 65241 40835 65307 40838
rect 65742 40836 65748 40838
rect 65812 40836 65818 40900
rect 65241 38722 65307 38725
rect 65926 38722 65932 38724
rect 65241 38720 65932 38722
rect 65241 38664 65246 38720
rect 65302 38664 65932 38720
rect 65241 38662 65932 38664
rect 65241 38659 65307 38662
rect 65926 38660 65932 38662
rect 65996 38660 66002 38724
rect 964 34592 75028 34616
rect 964 34588 4740 34592
rect 964 34532 2044 34588
rect 2100 34532 4740 34588
rect 964 34528 4740 34532
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34588 10740 34592
rect 5284 34532 5540 34588
rect 5596 34532 8430 34588
rect 8486 34532 10740 34588
rect 5284 34528 10740 34532
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34588 16740 34592
rect 11284 34532 11320 34588
rect 11376 34532 14210 34588
rect 14266 34532 16740 34588
rect 11284 34528 16740 34532
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34588 17140 34592
rect 17124 34528 17140 34532
rect 17204 34528 17220 34592
rect 17284 34588 22740 34592
rect 17284 34532 19990 34588
rect 20046 34532 22740 34588
rect 17284 34528 22740 34532
rect 22804 34528 22820 34592
rect 22884 34588 22900 34592
rect 22884 34528 22900 34532
rect 22964 34528 22980 34592
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34588 28740 34592
rect 23284 34532 25770 34588
rect 25826 34532 28660 34588
rect 28716 34532 28740 34588
rect 23284 34528 28740 34532
rect 28804 34528 28820 34592
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34588 34740 34592
rect 29284 34532 31550 34588
rect 31606 34532 34440 34588
rect 34496 34532 34740 34588
rect 29284 34528 34740 34532
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34588 40740 34592
rect 35284 34532 37330 34588
rect 37386 34532 40220 34588
rect 40276 34532 40740 34588
rect 35284 34528 40740 34532
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34588 46740 34592
rect 41284 34532 43110 34588
rect 43166 34532 46000 34588
rect 46056 34532 46740 34588
rect 41284 34528 46740 34532
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34588 52740 34592
rect 47284 34532 49008 34588
rect 49064 34532 52237 34588
rect 52293 34532 52740 34588
rect 47284 34528 52740 34532
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34588 58740 34592
rect 53284 34532 53638 34588
rect 53694 34532 53806 34588
rect 53862 34532 54550 34588
rect 54606 34532 54940 34588
rect 54996 34532 55656 34588
rect 55712 34532 56234 34588
rect 56290 34532 56679 34588
rect 56735 34532 56983 34588
rect 57039 34532 57825 34588
rect 57881 34532 58465 34588
rect 58521 34532 58740 34588
rect 53284 34528 58740 34532
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34588 59060 34592
rect 59044 34532 59048 34588
rect 59044 34528 59060 34532
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34588 64740 34592
rect 59284 34532 60326 34588
rect 60382 34532 60484 34588
rect 60540 34532 62528 34588
rect 62584 34532 62608 34588
rect 62664 34532 64740 34588
rect 59284 34528 64740 34532
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34588 75028 34592
rect 71284 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 75028 34588
rect 71284 34528 75028 34532
rect 964 34512 75028 34528
rect 964 34508 4740 34512
rect 964 34452 2044 34508
rect 2100 34452 4740 34508
rect 964 34448 4740 34452
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34508 10740 34512
rect 5284 34452 5540 34508
rect 5596 34452 8430 34508
rect 8486 34452 10740 34508
rect 5284 34448 10740 34452
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34508 16740 34512
rect 11284 34452 11320 34508
rect 11376 34452 14210 34508
rect 14266 34452 16740 34508
rect 11284 34448 16740 34452
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34508 17140 34512
rect 17124 34448 17140 34452
rect 17204 34448 17220 34512
rect 17284 34508 22740 34512
rect 17284 34452 19990 34508
rect 20046 34452 22740 34508
rect 17284 34448 22740 34452
rect 22804 34448 22820 34512
rect 22884 34508 22900 34512
rect 22884 34448 22900 34452
rect 22964 34448 22980 34512
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34508 28740 34512
rect 23284 34452 25770 34508
rect 25826 34452 28660 34508
rect 28716 34452 28740 34508
rect 23284 34448 28740 34452
rect 28804 34448 28820 34512
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34508 34740 34512
rect 29284 34452 31550 34508
rect 31606 34452 34440 34508
rect 34496 34452 34740 34508
rect 29284 34448 34740 34452
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34508 40740 34512
rect 35284 34452 37330 34508
rect 37386 34452 40220 34508
rect 40276 34452 40740 34508
rect 35284 34448 40740 34452
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34508 46740 34512
rect 41284 34452 43110 34508
rect 43166 34452 46000 34508
rect 46056 34452 46740 34508
rect 41284 34448 46740 34452
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34508 52740 34512
rect 47284 34452 49008 34508
rect 49064 34452 52237 34508
rect 52293 34452 52740 34508
rect 47284 34448 52740 34452
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34508 58740 34512
rect 53284 34452 53638 34508
rect 53694 34452 53806 34508
rect 53862 34452 54550 34508
rect 54606 34452 54940 34508
rect 54996 34452 55656 34508
rect 55712 34452 56234 34508
rect 56290 34452 56679 34508
rect 56735 34452 56983 34508
rect 57039 34452 57825 34508
rect 57881 34452 58465 34508
rect 58521 34452 58740 34508
rect 53284 34448 58740 34452
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34508 59060 34512
rect 59044 34452 59048 34508
rect 59044 34448 59060 34452
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34508 64740 34512
rect 59284 34452 60326 34508
rect 60382 34452 60484 34508
rect 60540 34452 62528 34508
rect 62584 34452 62608 34508
rect 62664 34452 64740 34508
rect 59284 34448 64740 34452
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34508 75028 34512
rect 71284 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 75028 34508
rect 71284 34448 75028 34452
rect 964 34432 75028 34448
rect 964 34428 4740 34432
rect 964 34372 2044 34428
rect 2100 34372 4740 34428
rect 964 34368 4740 34372
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34428 10740 34432
rect 5284 34372 5540 34428
rect 5596 34372 8430 34428
rect 8486 34372 10740 34428
rect 5284 34368 10740 34372
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34428 16740 34432
rect 11284 34372 11320 34428
rect 11376 34372 14210 34428
rect 14266 34372 16740 34428
rect 11284 34368 16740 34372
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34428 17140 34432
rect 17124 34368 17140 34372
rect 17204 34368 17220 34432
rect 17284 34428 22740 34432
rect 17284 34372 19990 34428
rect 20046 34372 22740 34428
rect 17284 34368 22740 34372
rect 22804 34368 22820 34432
rect 22884 34428 22900 34432
rect 22884 34368 22900 34372
rect 22964 34368 22980 34432
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34428 28740 34432
rect 23284 34372 25770 34428
rect 25826 34372 28660 34428
rect 28716 34372 28740 34428
rect 23284 34368 28740 34372
rect 28804 34368 28820 34432
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34428 34740 34432
rect 29284 34372 31550 34428
rect 31606 34372 34440 34428
rect 34496 34372 34740 34428
rect 29284 34368 34740 34372
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34428 40740 34432
rect 35284 34372 37330 34428
rect 37386 34372 40220 34428
rect 40276 34372 40740 34428
rect 35284 34368 40740 34372
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34428 46740 34432
rect 41284 34372 43110 34428
rect 43166 34372 46000 34428
rect 46056 34372 46740 34428
rect 41284 34368 46740 34372
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34428 52740 34432
rect 47284 34372 49008 34428
rect 49064 34372 52237 34428
rect 52293 34372 52740 34428
rect 47284 34368 52740 34372
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34428 58740 34432
rect 53284 34372 53638 34428
rect 53694 34372 53806 34428
rect 53862 34372 54550 34428
rect 54606 34372 54940 34428
rect 54996 34372 55656 34428
rect 55712 34372 56234 34428
rect 56290 34372 56679 34428
rect 56735 34372 56983 34428
rect 57039 34372 57825 34428
rect 57881 34372 58465 34428
rect 58521 34372 58740 34428
rect 53284 34368 58740 34372
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34428 59060 34432
rect 59044 34372 59048 34428
rect 59044 34368 59060 34372
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34428 64740 34432
rect 59284 34372 60326 34428
rect 60382 34372 60484 34428
rect 60540 34372 62528 34428
rect 62584 34372 62608 34428
rect 62664 34372 64740 34428
rect 59284 34368 64740 34372
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34428 75028 34432
rect 71284 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 75028 34428
rect 71284 34368 75028 34372
rect 964 34352 75028 34368
rect 964 34348 4740 34352
rect 964 34292 2044 34348
rect 2100 34292 4740 34348
rect 964 34288 4740 34292
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34348 10740 34352
rect 5284 34292 5540 34348
rect 5596 34292 8430 34348
rect 8486 34292 10740 34348
rect 5284 34288 10740 34292
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34348 16740 34352
rect 11284 34292 11320 34348
rect 11376 34292 14210 34348
rect 14266 34292 16740 34348
rect 11284 34288 16740 34292
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34348 17140 34352
rect 17124 34288 17140 34292
rect 17204 34288 17220 34352
rect 17284 34348 22740 34352
rect 17284 34292 19990 34348
rect 20046 34292 22740 34348
rect 17284 34288 22740 34292
rect 22804 34288 22820 34352
rect 22884 34348 22900 34352
rect 22884 34288 22900 34292
rect 22964 34288 22980 34352
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34348 28740 34352
rect 23284 34292 25770 34348
rect 25826 34292 28660 34348
rect 28716 34292 28740 34348
rect 23284 34288 28740 34292
rect 28804 34288 28820 34352
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34348 34740 34352
rect 29284 34292 31550 34348
rect 31606 34292 34440 34348
rect 34496 34292 34740 34348
rect 29284 34288 34740 34292
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34348 40740 34352
rect 35284 34292 37330 34348
rect 37386 34292 40220 34348
rect 40276 34292 40740 34348
rect 35284 34288 40740 34292
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34348 46740 34352
rect 41284 34292 43110 34348
rect 43166 34292 46000 34348
rect 46056 34292 46740 34348
rect 41284 34288 46740 34292
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34348 52740 34352
rect 47284 34292 49008 34348
rect 49064 34292 52237 34348
rect 52293 34292 52740 34348
rect 47284 34288 52740 34292
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34348 58740 34352
rect 53284 34292 53638 34348
rect 53694 34292 53806 34348
rect 53862 34292 54550 34348
rect 54606 34292 54940 34348
rect 54996 34292 55656 34348
rect 55712 34292 56234 34348
rect 56290 34292 56679 34348
rect 56735 34292 56983 34348
rect 57039 34292 57825 34348
rect 57881 34292 58465 34348
rect 58521 34292 58740 34348
rect 53284 34288 58740 34292
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34348 59060 34352
rect 59044 34292 59048 34348
rect 59044 34288 59060 34292
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34348 64740 34352
rect 59284 34292 60326 34348
rect 60382 34292 60484 34348
rect 60540 34292 62528 34348
rect 62584 34292 62608 34348
rect 62664 34292 64740 34348
rect 59284 34288 64740 34292
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34348 75028 34352
rect 71284 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 75028 34348
rect 71284 34288 75028 34292
rect 964 34264 75028 34288
rect 65609 33282 65675 33285
rect 68502 33282 68508 33284
rect 65609 33280 68508 33282
rect 65609 33224 65614 33280
rect 65670 33224 68508 33280
rect 65609 33222 68508 33224
rect 65609 33219 65675 33222
rect 68502 33220 68508 33222
rect 68572 33220 68578 33284
rect 964 32240 75028 32264
rect 964 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32236 2220 32240
rect 2284 32236 7740 32240
rect 2320 32180 5393 32236
rect 5449 32180 7740 32236
rect 2204 32176 2220 32180
rect 2284 32176 7740 32180
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32236 13740 32240
rect 8339 32180 11173 32236
rect 11229 32180 13740 32236
rect 8284 32176 13740 32180
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32176 14220 32240
rect 14284 32236 19740 32240
rect 14284 32180 16953 32236
rect 17009 32180 19740 32236
rect 14284 32176 19740 32180
rect 19804 32176 19820 32240
rect 19884 32236 19900 32240
rect 19899 32180 19900 32236
rect 19884 32176 19900 32180
rect 19964 32176 19980 32240
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32236 25740 32240
rect 20284 32180 22733 32236
rect 22789 32180 25623 32236
rect 25679 32180 25740 32236
rect 20284 32176 25740 32180
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32236 31740 32240
rect 26284 32180 28513 32236
rect 28569 32180 31403 32236
rect 31459 32180 31740 32236
rect 26284 32176 31740 32180
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32236 37740 32240
rect 32284 32180 34293 32236
rect 34349 32180 37183 32236
rect 37239 32180 37740 32236
rect 32284 32176 37740 32180
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32236 43740 32240
rect 38284 32180 40073 32236
rect 40129 32180 42963 32236
rect 43019 32180 43740 32236
rect 38284 32176 43740 32180
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32236 49740 32240
rect 44284 32180 45853 32236
rect 45909 32180 48800 32236
rect 48856 32180 49662 32236
rect 49718 32180 49740 32236
rect 44284 32176 49740 32180
rect 49804 32176 49820 32240
rect 49884 32176 49900 32240
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32236 55740 32240
rect 50284 32180 52956 32236
rect 53012 32180 53114 32236
rect 53170 32180 53470 32236
rect 53526 32180 54788 32236
rect 54844 32180 55381 32236
rect 55437 32180 55740 32236
rect 50284 32176 55740 32180
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32236 61740 32240
rect 56284 32180 56527 32236
rect 56583 32180 57963 32236
rect 58019 32180 58043 32236
rect 58099 32180 59206 32236
rect 59262 32180 59364 32236
rect 59420 32180 59672 32236
rect 59728 32180 59818 32236
rect 59874 32180 59954 32236
rect 60010 32180 60034 32236
rect 60090 32180 61740 32236
rect 56284 32176 61740 32180
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32236 67740 32240
rect 62284 32180 62326 32236
rect 62382 32180 62406 32236
rect 62462 32180 67740 32236
rect 62284 32176 67740 32180
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32236 73740 32240
rect 68284 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 73740 32236
rect 68284 32176 73740 32180
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 75028 32240
rect 964 32160 75028 32176
rect 964 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32156 2220 32160
rect 2284 32156 7740 32160
rect 2320 32100 5393 32156
rect 5449 32100 7740 32156
rect 2204 32096 2220 32100
rect 2284 32096 7740 32100
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32156 13740 32160
rect 8339 32100 11173 32156
rect 11229 32100 13740 32156
rect 8284 32096 13740 32100
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32096 14220 32160
rect 14284 32156 19740 32160
rect 14284 32100 16953 32156
rect 17009 32100 19740 32156
rect 14284 32096 19740 32100
rect 19804 32096 19820 32160
rect 19884 32156 19900 32160
rect 19899 32100 19900 32156
rect 19884 32096 19900 32100
rect 19964 32096 19980 32160
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32156 25740 32160
rect 20284 32100 22733 32156
rect 22789 32100 25623 32156
rect 25679 32100 25740 32156
rect 20284 32096 25740 32100
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32156 31740 32160
rect 26284 32100 28513 32156
rect 28569 32100 31403 32156
rect 31459 32100 31740 32156
rect 26284 32096 31740 32100
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32156 37740 32160
rect 32284 32100 34293 32156
rect 34349 32100 37183 32156
rect 37239 32100 37740 32156
rect 32284 32096 37740 32100
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32156 43740 32160
rect 38284 32100 40073 32156
rect 40129 32100 42963 32156
rect 43019 32100 43740 32156
rect 38284 32096 43740 32100
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32156 49740 32160
rect 44284 32100 45853 32156
rect 45909 32100 48800 32156
rect 48856 32100 49662 32156
rect 49718 32100 49740 32156
rect 44284 32096 49740 32100
rect 49804 32096 49820 32160
rect 49884 32096 49900 32160
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32156 55740 32160
rect 50284 32100 52956 32156
rect 53012 32100 53114 32156
rect 53170 32100 53470 32156
rect 53526 32100 54788 32156
rect 54844 32100 55381 32156
rect 55437 32100 55740 32156
rect 50284 32096 55740 32100
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32156 61740 32160
rect 56284 32100 56527 32156
rect 56583 32100 57963 32156
rect 58019 32100 58043 32156
rect 58099 32100 59206 32156
rect 59262 32100 59364 32156
rect 59420 32100 59672 32156
rect 59728 32100 59818 32156
rect 59874 32100 59954 32156
rect 60010 32100 60034 32156
rect 60090 32100 61740 32156
rect 56284 32096 61740 32100
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32156 67740 32160
rect 62284 32100 62326 32156
rect 62382 32100 62406 32156
rect 62462 32100 67740 32156
rect 62284 32096 67740 32100
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32156 73740 32160
rect 68284 32100 71864 32156
rect 71920 32100 71944 32156
rect 72000 32100 72024 32156
rect 72080 32100 72104 32156
rect 72160 32100 73740 32156
rect 68284 32096 73740 32100
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 75028 32160
rect 964 32080 75028 32096
rect 964 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32076 2220 32080
rect 2284 32076 7740 32080
rect 2320 32020 5393 32076
rect 5449 32020 7740 32076
rect 2204 32016 2220 32020
rect 2284 32016 7740 32020
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32076 13740 32080
rect 8339 32020 11173 32076
rect 11229 32020 13740 32076
rect 8284 32016 13740 32020
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32016 14220 32080
rect 14284 32076 19740 32080
rect 14284 32020 16953 32076
rect 17009 32020 19740 32076
rect 14284 32016 19740 32020
rect 19804 32016 19820 32080
rect 19884 32076 19900 32080
rect 19899 32020 19900 32076
rect 19884 32016 19900 32020
rect 19964 32016 19980 32080
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32076 25740 32080
rect 20284 32020 22733 32076
rect 22789 32020 25623 32076
rect 25679 32020 25740 32076
rect 20284 32016 25740 32020
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32076 31740 32080
rect 26284 32020 28513 32076
rect 28569 32020 31403 32076
rect 31459 32020 31740 32076
rect 26284 32016 31740 32020
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32076 37740 32080
rect 32284 32020 34293 32076
rect 34349 32020 37183 32076
rect 37239 32020 37740 32076
rect 32284 32016 37740 32020
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32076 43740 32080
rect 38284 32020 40073 32076
rect 40129 32020 42963 32076
rect 43019 32020 43740 32076
rect 38284 32016 43740 32020
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32076 49740 32080
rect 44284 32020 45853 32076
rect 45909 32020 48800 32076
rect 48856 32020 49662 32076
rect 49718 32020 49740 32076
rect 44284 32016 49740 32020
rect 49804 32016 49820 32080
rect 49884 32016 49900 32080
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32076 55740 32080
rect 50284 32020 52956 32076
rect 53012 32020 53114 32076
rect 53170 32020 53470 32076
rect 53526 32020 54788 32076
rect 54844 32020 55381 32076
rect 55437 32020 55740 32076
rect 50284 32016 55740 32020
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32076 61740 32080
rect 56284 32020 56527 32076
rect 56583 32020 57963 32076
rect 58019 32020 58043 32076
rect 58099 32020 59206 32076
rect 59262 32020 59364 32076
rect 59420 32020 59672 32076
rect 59728 32020 59818 32076
rect 59874 32020 59954 32076
rect 60010 32020 60034 32076
rect 60090 32020 61740 32076
rect 56284 32016 61740 32020
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32076 67740 32080
rect 62284 32020 62326 32076
rect 62382 32020 62406 32076
rect 62462 32020 67740 32076
rect 62284 32016 67740 32020
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32076 73740 32080
rect 68284 32020 71864 32076
rect 71920 32020 71944 32076
rect 72000 32020 72024 32076
rect 72080 32020 72104 32076
rect 72160 32020 73740 32076
rect 68284 32016 73740 32020
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 75028 32080
rect 964 32000 75028 32016
rect 964 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31996 2220 32000
rect 2284 31996 7740 32000
rect 2320 31940 5393 31996
rect 5449 31940 7740 31996
rect 2204 31936 2220 31940
rect 2284 31936 7740 31940
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31996 13740 32000
rect 8339 31940 11173 31996
rect 11229 31940 13740 31996
rect 8284 31936 13740 31940
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31936 14220 32000
rect 14284 31996 19740 32000
rect 14284 31940 16953 31996
rect 17009 31940 19740 31996
rect 14284 31936 19740 31940
rect 19804 31936 19820 32000
rect 19884 31996 19900 32000
rect 19899 31940 19900 31996
rect 19884 31936 19900 31940
rect 19964 31936 19980 32000
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31996 25740 32000
rect 20284 31940 22733 31996
rect 22789 31940 25623 31996
rect 25679 31940 25740 31996
rect 20284 31936 25740 31940
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31996 31740 32000
rect 26284 31940 28513 31996
rect 28569 31940 31403 31996
rect 31459 31940 31740 31996
rect 26284 31936 31740 31940
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31996 37740 32000
rect 32284 31940 34293 31996
rect 34349 31940 37183 31996
rect 37239 31940 37740 31996
rect 32284 31936 37740 31940
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31996 43740 32000
rect 38284 31940 40073 31996
rect 40129 31940 42963 31996
rect 43019 31940 43740 31996
rect 38284 31936 43740 31940
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31996 49740 32000
rect 44284 31940 45853 31996
rect 45909 31940 48800 31996
rect 48856 31940 49662 31996
rect 49718 31940 49740 31996
rect 44284 31936 49740 31940
rect 49804 31936 49820 32000
rect 49884 31936 49900 32000
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31996 55740 32000
rect 50284 31940 52956 31996
rect 53012 31940 53114 31996
rect 53170 31940 53470 31996
rect 53526 31940 54788 31996
rect 54844 31940 55381 31996
rect 55437 31940 55740 31996
rect 50284 31936 55740 31940
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31996 61740 32000
rect 56284 31940 56527 31996
rect 56583 31940 57963 31996
rect 58019 31940 58043 31996
rect 58099 31940 59206 31996
rect 59262 31940 59364 31996
rect 59420 31940 59672 31996
rect 59728 31940 59818 31996
rect 59874 31940 59954 31996
rect 60010 31940 60034 31996
rect 60090 31940 61740 31996
rect 56284 31936 61740 31940
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31996 67740 32000
rect 62284 31940 62326 31996
rect 62382 31940 62406 31996
rect 62462 31940 67740 31996
rect 62284 31936 67740 31940
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31996 73740 32000
rect 68284 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 73740 31996
rect 68284 31936 73740 31940
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 75028 32000
rect 964 31912 75028 31936
rect 964 24592 75028 24616
rect 964 24588 4740 24592
rect 964 24532 2044 24588
rect 2100 24532 4740 24588
rect 964 24528 4740 24532
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24588 10740 24592
rect 5284 24532 5540 24588
rect 5596 24532 8430 24588
rect 8486 24532 10740 24588
rect 5284 24528 10740 24532
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24588 16740 24592
rect 11284 24532 11320 24588
rect 11376 24532 14210 24588
rect 14266 24532 16740 24588
rect 11284 24528 16740 24532
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24588 17140 24592
rect 17124 24528 17140 24532
rect 17204 24528 17220 24592
rect 17284 24588 22740 24592
rect 17284 24532 19990 24588
rect 20046 24532 22740 24588
rect 17284 24528 22740 24532
rect 22804 24528 22820 24592
rect 22884 24588 22900 24592
rect 22884 24528 22900 24532
rect 22964 24528 22980 24592
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24588 28740 24592
rect 23284 24532 25770 24588
rect 25826 24532 28660 24588
rect 28716 24532 28740 24588
rect 23284 24528 28740 24532
rect 28804 24528 28820 24592
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24588 34740 24592
rect 29284 24532 31550 24588
rect 31606 24532 34440 24588
rect 34496 24532 34740 24588
rect 29284 24528 34740 24532
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24588 40740 24592
rect 35284 24532 37330 24588
rect 37386 24532 40220 24588
rect 40276 24532 40740 24588
rect 35284 24528 40740 24532
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24588 46740 24592
rect 41284 24532 43110 24588
rect 43166 24532 46000 24588
rect 46056 24532 46740 24588
rect 41284 24528 46740 24532
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24588 52740 24592
rect 47284 24532 49008 24588
rect 49064 24532 52237 24588
rect 52293 24532 52740 24588
rect 47284 24528 52740 24532
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24588 58740 24592
rect 53284 24532 53638 24588
rect 53694 24532 53806 24588
rect 53862 24532 54550 24588
rect 54606 24532 54940 24588
rect 54996 24532 55656 24588
rect 55712 24532 56234 24588
rect 56290 24532 56679 24588
rect 56735 24532 56983 24588
rect 57039 24532 57825 24588
rect 57881 24532 58465 24588
rect 58521 24532 58740 24588
rect 53284 24528 58740 24532
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24588 59060 24592
rect 59044 24532 59048 24588
rect 59044 24528 59060 24532
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24588 64740 24592
rect 59284 24532 60326 24588
rect 60382 24532 60484 24588
rect 60540 24532 62528 24588
rect 62584 24532 62608 24588
rect 62664 24532 64740 24588
rect 59284 24528 64740 24532
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24588 75028 24592
rect 71284 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 75028 24588
rect 71284 24528 75028 24532
rect 964 24512 75028 24528
rect 964 24508 4740 24512
rect 964 24452 2044 24508
rect 2100 24452 4740 24508
rect 964 24448 4740 24452
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24508 10740 24512
rect 5284 24452 5540 24508
rect 5596 24452 8430 24508
rect 8486 24452 10740 24508
rect 5284 24448 10740 24452
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24508 16740 24512
rect 11284 24452 11320 24508
rect 11376 24452 14210 24508
rect 14266 24452 16740 24508
rect 11284 24448 16740 24452
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24508 17140 24512
rect 17124 24448 17140 24452
rect 17204 24448 17220 24512
rect 17284 24508 22740 24512
rect 17284 24452 19990 24508
rect 20046 24452 22740 24508
rect 17284 24448 22740 24452
rect 22804 24448 22820 24512
rect 22884 24508 22900 24512
rect 22884 24448 22900 24452
rect 22964 24448 22980 24512
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24508 28740 24512
rect 23284 24452 25770 24508
rect 25826 24452 28660 24508
rect 28716 24452 28740 24508
rect 23284 24448 28740 24452
rect 28804 24448 28820 24512
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24508 34740 24512
rect 29284 24452 31550 24508
rect 31606 24452 34440 24508
rect 34496 24452 34740 24508
rect 29284 24448 34740 24452
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24508 40740 24512
rect 35284 24452 37330 24508
rect 37386 24452 40220 24508
rect 40276 24452 40740 24508
rect 35284 24448 40740 24452
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24508 46740 24512
rect 41284 24452 43110 24508
rect 43166 24452 46000 24508
rect 46056 24452 46740 24508
rect 41284 24448 46740 24452
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24508 52740 24512
rect 47284 24452 49008 24508
rect 49064 24452 52237 24508
rect 52293 24452 52740 24508
rect 47284 24448 52740 24452
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24508 58740 24512
rect 53284 24452 53638 24508
rect 53694 24452 53806 24508
rect 53862 24452 54550 24508
rect 54606 24452 54940 24508
rect 54996 24452 55656 24508
rect 55712 24452 56234 24508
rect 56290 24452 56679 24508
rect 56735 24452 56983 24508
rect 57039 24452 57825 24508
rect 57881 24452 58465 24508
rect 58521 24452 58740 24508
rect 53284 24448 58740 24452
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24508 59060 24512
rect 59044 24452 59048 24508
rect 59044 24448 59060 24452
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24508 64740 24512
rect 59284 24452 60326 24508
rect 60382 24452 60484 24508
rect 60540 24452 62528 24508
rect 62584 24452 62608 24508
rect 62664 24452 64740 24508
rect 59284 24448 64740 24452
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24508 75028 24512
rect 71284 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 75028 24508
rect 71284 24448 75028 24452
rect 964 24432 75028 24448
rect 964 24428 4740 24432
rect 964 24372 2044 24428
rect 2100 24372 4740 24428
rect 964 24368 4740 24372
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24428 10740 24432
rect 5284 24372 5540 24428
rect 5596 24372 8430 24428
rect 8486 24372 10740 24428
rect 5284 24368 10740 24372
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24428 16740 24432
rect 11284 24372 11320 24428
rect 11376 24372 14210 24428
rect 14266 24372 16740 24428
rect 11284 24368 16740 24372
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24428 17140 24432
rect 17124 24368 17140 24372
rect 17204 24368 17220 24432
rect 17284 24428 22740 24432
rect 17284 24372 19990 24428
rect 20046 24372 22740 24428
rect 17284 24368 22740 24372
rect 22804 24368 22820 24432
rect 22884 24428 22900 24432
rect 22884 24368 22900 24372
rect 22964 24368 22980 24432
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24428 28740 24432
rect 23284 24372 25770 24428
rect 25826 24372 28660 24428
rect 28716 24372 28740 24428
rect 23284 24368 28740 24372
rect 28804 24368 28820 24432
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24428 34740 24432
rect 29284 24372 31550 24428
rect 31606 24372 34440 24428
rect 34496 24372 34740 24428
rect 29284 24368 34740 24372
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24428 40740 24432
rect 35284 24372 37330 24428
rect 37386 24372 40220 24428
rect 40276 24372 40740 24428
rect 35284 24368 40740 24372
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24428 46740 24432
rect 41284 24372 43110 24428
rect 43166 24372 46000 24428
rect 46056 24372 46740 24428
rect 41284 24368 46740 24372
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24428 52740 24432
rect 47284 24372 49008 24428
rect 49064 24372 52237 24428
rect 52293 24372 52740 24428
rect 47284 24368 52740 24372
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24428 58740 24432
rect 53284 24372 53638 24428
rect 53694 24372 53806 24428
rect 53862 24372 54550 24428
rect 54606 24372 54940 24428
rect 54996 24372 55656 24428
rect 55712 24372 56234 24428
rect 56290 24372 56679 24428
rect 56735 24372 56983 24428
rect 57039 24372 57825 24428
rect 57881 24372 58465 24428
rect 58521 24372 58740 24428
rect 53284 24368 58740 24372
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24428 59060 24432
rect 59044 24372 59048 24428
rect 59044 24368 59060 24372
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24428 64740 24432
rect 59284 24372 60326 24428
rect 60382 24372 60484 24428
rect 60540 24372 62528 24428
rect 62584 24372 62608 24428
rect 62664 24372 64740 24428
rect 59284 24368 64740 24372
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24428 75028 24432
rect 71284 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 75028 24428
rect 71284 24368 75028 24372
rect 964 24352 75028 24368
rect 964 24348 4740 24352
rect 964 24292 2044 24348
rect 2100 24292 4740 24348
rect 964 24288 4740 24292
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24348 10740 24352
rect 5284 24292 5540 24348
rect 5596 24292 8430 24348
rect 8486 24292 10740 24348
rect 5284 24288 10740 24292
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24348 16740 24352
rect 11284 24292 11320 24348
rect 11376 24292 14210 24348
rect 14266 24292 16740 24348
rect 11284 24288 16740 24292
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24348 17140 24352
rect 17124 24288 17140 24292
rect 17204 24288 17220 24352
rect 17284 24348 22740 24352
rect 17284 24292 19990 24348
rect 20046 24292 22740 24348
rect 17284 24288 22740 24292
rect 22804 24288 22820 24352
rect 22884 24348 22900 24352
rect 22884 24288 22900 24292
rect 22964 24288 22980 24352
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24348 28740 24352
rect 23284 24292 25770 24348
rect 25826 24292 28660 24348
rect 28716 24292 28740 24348
rect 23284 24288 28740 24292
rect 28804 24288 28820 24352
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24348 34740 24352
rect 29284 24292 31550 24348
rect 31606 24292 34440 24348
rect 34496 24292 34740 24348
rect 29284 24288 34740 24292
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24348 40740 24352
rect 35284 24292 37330 24348
rect 37386 24292 40220 24348
rect 40276 24292 40740 24348
rect 35284 24288 40740 24292
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24348 46740 24352
rect 41284 24292 43110 24348
rect 43166 24292 46000 24348
rect 46056 24292 46740 24348
rect 41284 24288 46740 24292
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24348 52740 24352
rect 47284 24292 49008 24348
rect 49064 24292 52237 24348
rect 52293 24292 52740 24348
rect 47284 24288 52740 24292
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24348 58740 24352
rect 53284 24292 53638 24348
rect 53694 24292 53806 24348
rect 53862 24292 54550 24348
rect 54606 24292 54940 24348
rect 54996 24292 55656 24348
rect 55712 24292 56234 24348
rect 56290 24292 56679 24348
rect 56735 24292 56983 24348
rect 57039 24292 57825 24348
rect 57881 24292 58465 24348
rect 58521 24292 58740 24348
rect 53284 24288 58740 24292
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24348 59060 24352
rect 59044 24292 59048 24348
rect 59044 24288 59060 24292
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24348 64740 24352
rect 59284 24292 60326 24348
rect 60382 24292 60484 24348
rect 60540 24292 62528 24348
rect 62584 24292 62608 24348
rect 62664 24292 64740 24348
rect 59284 24288 64740 24292
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24348 75028 24352
rect 71284 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 75028 24348
rect 71284 24288 75028 24292
rect 964 24264 75028 24288
rect 66989 23898 67055 23901
rect 66854 23896 67055 23898
rect 66854 23840 66994 23896
rect 67050 23840 67055 23896
rect 66854 23838 67055 23840
rect 66345 23492 66411 23493
rect 66529 23492 66595 23493
rect 66294 23490 66300 23492
rect 66254 23430 66300 23490
rect 66364 23488 66411 23492
rect 66406 23432 66411 23488
rect 66294 23428 66300 23430
rect 66364 23428 66411 23432
rect 66478 23428 66484 23492
rect 66548 23490 66595 23492
rect 66548 23488 66640 23490
rect 66590 23432 66640 23488
rect 66548 23430 66640 23432
rect 66548 23428 66595 23430
rect 66345 23427 66411 23428
rect 66529 23427 66595 23428
rect 66345 23354 66411 23357
rect 66854 23354 66914 23838
rect 66989 23835 67055 23838
rect 66345 23352 66914 23354
rect 66345 23296 66350 23352
rect 66406 23296 66914 23352
rect 66345 23294 66914 23296
rect 66345 23291 66411 23294
rect 964 22240 75028 22264
rect 964 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22236 2220 22240
rect 2284 22236 7740 22240
rect 2320 22180 5393 22236
rect 5449 22180 7740 22236
rect 2204 22176 2220 22180
rect 2284 22176 7740 22180
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22236 13740 22240
rect 8339 22180 11173 22236
rect 11229 22180 13740 22236
rect 8284 22176 13740 22180
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22176 14220 22240
rect 14284 22236 19740 22240
rect 14284 22180 16953 22236
rect 17009 22180 19740 22236
rect 14284 22176 19740 22180
rect 19804 22176 19820 22240
rect 19884 22236 19900 22240
rect 19899 22180 19900 22236
rect 19884 22176 19900 22180
rect 19964 22176 19980 22240
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22236 25740 22240
rect 20284 22180 22733 22236
rect 22789 22180 25623 22236
rect 25679 22180 25740 22236
rect 20284 22176 25740 22180
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22236 31740 22240
rect 26284 22180 28513 22236
rect 28569 22180 31403 22236
rect 31459 22180 31740 22236
rect 26284 22176 31740 22180
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22236 37740 22240
rect 32284 22180 34293 22236
rect 34349 22180 37183 22236
rect 37239 22180 37740 22236
rect 32284 22176 37740 22180
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22236 43740 22240
rect 38284 22180 40073 22236
rect 40129 22180 42963 22236
rect 43019 22180 43740 22236
rect 38284 22176 43740 22180
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22236 49740 22240
rect 44284 22180 45853 22236
rect 45909 22180 48800 22236
rect 48856 22180 49662 22236
rect 49718 22180 49740 22236
rect 44284 22176 49740 22180
rect 49804 22176 49820 22240
rect 49884 22176 49900 22240
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22236 55740 22240
rect 50284 22180 52956 22236
rect 53012 22180 53114 22236
rect 53170 22180 53470 22236
rect 53526 22180 54788 22236
rect 54844 22180 55381 22236
rect 55437 22180 55740 22236
rect 50284 22176 55740 22180
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22236 61740 22240
rect 56284 22180 56527 22236
rect 56583 22180 57963 22236
rect 58019 22180 58043 22236
rect 58099 22180 59206 22236
rect 59262 22180 59364 22236
rect 59420 22180 59672 22236
rect 59728 22180 59818 22236
rect 59874 22180 59954 22236
rect 60010 22180 60034 22236
rect 60090 22180 61740 22236
rect 56284 22176 61740 22180
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22236 67740 22240
rect 62284 22180 62326 22236
rect 62382 22180 62406 22236
rect 62462 22180 67740 22236
rect 62284 22176 67740 22180
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22236 73740 22240
rect 68284 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 73740 22236
rect 68284 22176 73740 22180
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 75028 22240
rect 964 22160 75028 22176
rect 964 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22156 2220 22160
rect 2284 22156 7740 22160
rect 2320 22100 5393 22156
rect 5449 22100 7740 22156
rect 2204 22096 2220 22100
rect 2284 22096 7740 22100
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22156 13740 22160
rect 8339 22100 11173 22156
rect 11229 22100 13740 22156
rect 8284 22096 13740 22100
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22096 14220 22160
rect 14284 22156 19740 22160
rect 14284 22100 16953 22156
rect 17009 22100 19740 22156
rect 14284 22096 19740 22100
rect 19804 22096 19820 22160
rect 19884 22156 19900 22160
rect 19899 22100 19900 22156
rect 19884 22096 19900 22100
rect 19964 22096 19980 22160
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22156 25740 22160
rect 20284 22100 22733 22156
rect 22789 22100 25623 22156
rect 25679 22100 25740 22156
rect 20284 22096 25740 22100
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22156 31740 22160
rect 26284 22100 28513 22156
rect 28569 22100 31403 22156
rect 31459 22100 31740 22156
rect 26284 22096 31740 22100
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22156 37740 22160
rect 32284 22100 34293 22156
rect 34349 22100 37183 22156
rect 37239 22100 37740 22156
rect 32284 22096 37740 22100
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22156 43740 22160
rect 38284 22100 40073 22156
rect 40129 22100 42963 22156
rect 43019 22100 43740 22156
rect 38284 22096 43740 22100
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22156 49740 22160
rect 44284 22100 45853 22156
rect 45909 22100 48800 22156
rect 48856 22100 49662 22156
rect 49718 22100 49740 22156
rect 44284 22096 49740 22100
rect 49804 22096 49820 22160
rect 49884 22096 49900 22160
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22156 55740 22160
rect 50284 22100 52956 22156
rect 53012 22100 53114 22156
rect 53170 22100 53470 22156
rect 53526 22100 54788 22156
rect 54844 22100 55381 22156
rect 55437 22100 55740 22156
rect 50284 22096 55740 22100
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22156 61740 22160
rect 56284 22100 56527 22156
rect 56583 22100 57963 22156
rect 58019 22100 58043 22156
rect 58099 22100 59206 22156
rect 59262 22100 59364 22156
rect 59420 22100 59672 22156
rect 59728 22100 59818 22156
rect 59874 22100 59954 22156
rect 60010 22100 60034 22156
rect 60090 22100 61740 22156
rect 56284 22096 61740 22100
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22156 67740 22160
rect 62284 22100 62326 22156
rect 62382 22100 62406 22156
rect 62462 22100 67740 22156
rect 62284 22096 67740 22100
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22156 73740 22160
rect 68284 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 73740 22156
rect 68284 22096 73740 22100
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 75028 22160
rect 964 22080 75028 22096
rect 964 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22076 2220 22080
rect 2284 22076 7740 22080
rect 2320 22020 5393 22076
rect 5449 22020 7740 22076
rect 2204 22016 2220 22020
rect 2284 22016 7740 22020
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22076 13740 22080
rect 8339 22020 11173 22076
rect 11229 22020 13740 22076
rect 8284 22016 13740 22020
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22016 14220 22080
rect 14284 22076 19740 22080
rect 14284 22020 16953 22076
rect 17009 22020 19740 22076
rect 14284 22016 19740 22020
rect 19804 22016 19820 22080
rect 19884 22076 19900 22080
rect 19899 22020 19900 22076
rect 19884 22016 19900 22020
rect 19964 22016 19980 22080
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22076 25740 22080
rect 20284 22020 22733 22076
rect 22789 22020 25623 22076
rect 25679 22020 25740 22076
rect 20284 22016 25740 22020
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22076 31740 22080
rect 26284 22020 28513 22076
rect 28569 22020 31403 22076
rect 31459 22020 31740 22076
rect 26284 22016 31740 22020
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22076 37740 22080
rect 32284 22020 34293 22076
rect 34349 22020 37183 22076
rect 37239 22020 37740 22076
rect 32284 22016 37740 22020
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22076 43740 22080
rect 38284 22020 40073 22076
rect 40129 22020 42963 22076
rect 43019 22020 43740 22076
rect 38284 22016 43740 22020
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22076 49740 22080
rect 44284 22020 45853 22076
rect 45909 22020 48800 22076
rect 48856 22020 49662 22076
rect 49718 22020 49740 22076
rect 44284 22016 49740 22020
rect 49804 22016 49820 22080
rect 49884 22016 49900 22080
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22076 55740 22080
rect 50284 22020 52956 22076
rect 53012 22020 53114 22076
rect 53170 22020 53470 22076
rect 53526 22020 54788 22076
rect 54844 22020 55381 22076
rect 55437 22020 55740 22076
rect 50284 22016 55740 22020
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22076 61740 22080
rect 56284 22020 56527 22076
rect 56583 22020 57963 22076
rect 58019 22020 58043 22076
rect 58099 22020 59206 22076
rect 59262 22020 59364 22076
rect 59420 22020 59672 22076
rect 59728 22020 59818 22076
rect 59874 22020 59954 22076
rect 60010 22020 60034 22076
rect 60090 22020 61740 22076
rect 56284 22016 61740 22020
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22076 67740 22080
rect 62284 22020 62326 22076
rect 62382 22020 62406 22076
rect 62462 22020 67740 22076
rect 62284 22016 67740 22020
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22076 73740 22080
rect 68284 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 73740 22076
rect 68284 22016 73740 22020
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 75028 22080
rect 964 22000 75028 22016
rect 964 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21996 2220 22000
rect 2284 21996 7740 22000
rect 2320 21940 5393 21996
rect 5449 21940 7740 21996
rect 2204 21936 2220 21940
rect 2284 21936 7740 21940
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21996 13740 22000
rect 8339 21940 11173 21996
rect 11229 21940 13740 21996
rect 8284 21936 13740 21940
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21936 14220 22000
rect 14284 21996 19740 22000
rect 14284 21940 16953 21996
rect 17009 21940 19740 21996
rect 14284 21936 19740 21940
rect 19804 21936 19820 22000
rect 19884 21996 19900 22000
rect 19899 21940 19900 21996
rect 19884 21936 19900 21940
rect 19964 21936 19980 22000
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21996 25740 22000
rect 20284 21940 22733 21996
rect 22789 21940 25623 21996
rect 25679 21940 25740 21996
rect 20284 21936 25740 21940
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21996 31740 22000
rect 26284 21940 28513 21996
rect 28569 21940 31403 21996
rect 31459 21940 31740 21996
rect 26284 21936 31740 21940
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21996 37740 22000
rect 32284 21940 34293 21996
rect 34349 21940 37183 21996
rect 37239 21940 37740 21996
rect 32284 21936 37740 21940
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21996 43740 22000
rect 38284 21940 40073 21996
rect 40129 21940 42963 21996
rect 43019 21940 43740 21996
rect 38284 21936 43740 21940
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21996 49740 22000
rect 44284 21940 45853 21996
rect 45909 21940 48800 21996
rect 48856 21940 49662 21996
rect 49718 21940 49740 21996
rect 44284 21936 49740 21940
rect 49804 21936 49820 22000
rect 49884 21936 49900 22000
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21996 55740 22000
rect 50284 21940 52956 21996
rect 53012 21940 53114 21996
rect 53170 21940 53470 21996
rect 53526 21940 54788 21996
rect 54844 21940 55381 21996
rect 55437 21940 55740 21996
rect 50284 21936 55740 21940
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21996 61740 22000
rect 56284 21940 56527 21996
rect 56583 21940 57963 21996
rect 58019 21940 58043 21996
rect 58099 21940 59206 21996
rect 59262 21940 59364 21996
rect 59420 21940 59672 21996
rect 59728 21940 59818 21996
rect 59874 21940 59954 21996
rect 60010 21940 60034 21996
rect 60090 21940 61740 21996
rect 56284 21936 61740 21940
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21996 67740 22000
rect 62284 21940 62326 21996
rect 62382 21940 62406 21996
rect 62462 21940 67740 21996
rect 62284 21936 67740 21940
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21996 73740 22000
rect 68284 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 73740 21996
rect 68284 21936 73740 21940
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 75028 22000
rect 964 21912 75028 21936
rect 65517 19138 65583 19141
rect 66662 19138 66668 19140
rect 65517 19136 66668 19138
rect 65517 19080 65522 19136
rect 65578 19080 66668 19136
rect 65517 19078 66668 19080
rect 65517 19075 65583 19078
rect 66662 19076 66668 19078
rect 66732 19076 66738 19140
rect 62982 17852 62988 17916
rect 63052 17914 63058 17916
rect 63677 17914 63743 17917
rect 63052 17912 63743 17914
rect 63052 17856 63682 17912
rect 63738 17856 63743 17912
rect 63052 17854 63743 17856
rect 63052 17852 63058 17854
rect 63677 17851 63743 17854
rect 964 14592 75028 14616
rect 964 14588 4740 14592
rect 964 14532 2044 14588
rect 2100 14532 4740 14588
rect 964 14528 4740 14532
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14588 10740 14592
rect 5284 14532 5540 14588
rect 5596 14532 8430 14588
rect 8486 14532 10740 14588
rect 5284 14528 10740 14532
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14588 16740 14592
rect 11284 14532 11320 14588
rect 11376 14532 14210 14588
rect 14266 14532 16740 14588
rect 11284 14528 16740 14532
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14588 17140 14592
rect 17124 14528 17140 14532
rect 17204 14528 17220 14592
rect 17284 14588 22740 14592
rect 17284 14532 19990 14588
rect 20046 14532 22740 14588
rect 17284 14528 22740 14532
rect 22804 14528 22820 14592
rect 22884 14588 22900 14592
rect 22884 14528 22900 14532
rect 22964 14528 22980 14592
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14588 28740 14592
rect 23284 14532 25770 14588
rect 25826 14532 28660 14588
rect 28716 14532 28740 14588
rect 23284 14528 28740 14532
rect 28804 14528 28820 14592
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14588 34740 14592
rect 29284 14532 31550 14588
rect 31606 14532 34440 14588
rect 34496 14532 34740 14588
rect 29284 14528 34740 14532
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14588 40740 14592
rect 35284 14532 37330 14588
rect 37386 14532 40220 14588
rect 40276 14532 40740 14588
rect 35284 14528 40740 14532
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14588 46740 14592
rect 41284 14532 43110 14588
rect 43166 14532 46000 14588
rect 46056 14532 46740 14588
rect 41284 14528 46740 14532
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14588 52740 14592
rect 47284 14532 49008 14588
rect 49064 14532 52237 14588
rect 52293 14532 52740 14588
rect 47284 14528 52740 14532
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14588 58740 14592
rect 53284 14532 53638 14588
rect 53694 14532 53806 14588
rect 53862 14532 54550 14588
rect 54606 14532 54940 14588
rect 54996 14532 55656 14588
rect 55712 14532 56234 14588
rect 56290 14532 56679 14588
rect 56735 14532 56983 14588
rect 57039 14532 57825 14588
rect 57881 14532 58465 14588
rect 58521 14532 58740 14588
rect 53284 14528 58740 14532
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14588 59060 14592
rect 59044 14532 59048 14588
rect 59044 14528 59060 14532
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14588 64740 14592
rect 59284 14532 60326 14588
rect 60382 14532 60484 14588
rect 60540 14532 62528 14588
rect 62584 14532 62608 14588
rect 62664 14532 64740 14588
rect 59284 14528 64740 14532
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14588 75028 14592
rect 71284 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 75028 14588
rect 71284 14528 75028 14532
rect 964 14512 75028 14528
rect 964 14508 4740 14512
rect 964 14452 2044 14508
rect 2100 14452 4740 14508
rect 964 14448 4740 14452
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14508 10740 14512
rect 5284 14452 5540 14508
rect 5596 14452 8430 14508
rect 8486 14452 10740 14508
rect 5284 14448 10740 14452
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14508 16740 14512
rect 11284 14452 11320 14508
rect 11376 14452 14210 14508
rect 14266 14452 16740 14508
rect 11284 14448 16740 14452
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14508 17140 14512
rect 17124 14448 17140 14452
rect 17204 14448 17220 14512
rect 17284 14508 22740 14512
rect 17284 14452 19990 14508
rect 20046 14452 22740 14508
rect 17284 14448 22740 14452
rect 22804 14448 22820 14512
rect 22884 14508 22900 14512
rect 22884 14448 22900 14452
rect 22964 14448 22980 14512
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14508 28740 14512
rect 23284 14452 25770 14508
rect 25826 14452 28660 14508
rect 28716 14452 28740 14508
rect 23284 14448 28740 14452
rect 28804 14448 28820 14512
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14508 34740 14512
rect 29284 14452 31550 14508
rect 31606 14452 34440 14508
rect 34496 14452 34740 14508
rect 29284 14448 34740 14452
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14508 40740 14512
rect 35284 14452 37330 14508
rect 37386 14452 40220 14508
rect 40276 14452 40740 14508
rect 35284 14448 40740 14452
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14508 46740 14512
rect 41284 14452 43110 14508
rect 43166 14452 46000 14508
rect 46056 14452 46740 14508
rect 41284 14448 46740 14452
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14508 52740 14512
rect 47284 14452 49008 14508
rect 49064 14452 52237 14508
rect 52293 14452 52740 14508
rect 47284 14448 52740 14452
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14508 58740 14512
rect 53284 14452 53638 14508
rect 53694 14452 53806 14508
rect 53862 14452 54550 14508
rect 54606 14452 54940 14508
rect 54996 14452 55656 14508
rect 55712 14452 56234 14508
rect 56290 14452 56679 14508
rect 56735 14452 56983 14508
rect 57039 14452 57825 14508
rect 57881 14452 58465 14508
rect 58521 14452 58740 14508
rect 53284 14448 58740 14452
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14508 59060 14512
rect 59044 14452 59048 14508
rect 59044 14448 59060 14452
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14508 64740 14512
rect 59284 14452 60326 14508
rect 60382 14452 60484 14508
rect 60540 14452 62528 14508
rect 62584 14452 62608 14508
rect 62664 14452 64740 14508
rect 59284 14448 64740 14452
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14508 75028 14512
rect 71284 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 75028 14508
rect 71284 14448 75028 14452
rect 964 14432 75028 14448
rect 964 14428 4740 14432
rect 964 14372 2044 14428
rect 2100 14372 4740 14428
rect 964 14368 4740 14372
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14428 10740 14432
rect 5284 14372 5540 14428
rect 5596 14372 8430 14428
rect 8486 14372 10740 14428
rect 5284 14368 10740 14372
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14428 16740 14432
rect 11284 14372 11320 14428
rect 11376 14372 14210 14428
rect 14266 14372 16740 14428
rect 11284 14368 16740 14372
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14428 17140 14432
rect 17124 14368 17140 14372
rect 17204 14368 17220 14432
rect 17284 14428 22740 14432
rect 17284 14372 19990 14428
rect 20046 14372 22740 14428
rect 17284 14368 22740 14372
rect 22804 14368 22820 14432
rect 22884 14428 22900 14432
rect 22884 14368 22900 14372
rect 22964 14368 22980 14432
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14428 28740 14432
rect 23284 14372 25770 14428
rect 25826 14372 28660 14428
rect 28716 14372 28740 14428
rect 23284 14368 28740 14372
rect 28804 14368 28820 14432
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14428 34740 14432
rect 29284 14372 31550 14428
rect 31606 14372 34440 14428
rect 34496 14372 34740 14428
rect 29284 14368 34740 14372
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14428 40740 14432
rect 35284 14372 37330 14428
rect 37386 14372 40220 14428
rect 40276 14372 40740 14428
rect 35284 14368 40740 14372
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14428 46740 14432
rect 41284 14372 43110 14428
rect 43166 14372 46000 14428
rect 46056 14372 46740 14428
rect 41284 14368 46740 14372
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14428 52740 14432
rect 47284 14372 49008 14428
rect 49064 14372 52237 14428
rect 52293 14372 52740 14428
rect 47284 14368 52740 14372
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14428 58740 14432
rect 53284 14372 53638 14428
rect 53694 14372 53806 14428
rect 53862 14372 54550 14428
rect 54606 14372 54940 14428
rect 54996 14372 55656 14428
rect 55712 14372 56234 14428
rect 56290 14372 56679 14428
rect 56735 14372 56983 14428
rect 57039 14372 57825 14428
rect 57881 14372 58465 14428
rect 58521 14372 58740 14428
rect 53284 14368 58740 14372
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14428 59060 14432
rect 59044 14372 59048 14428
rect 59044 14368 59060 14372
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14428 64740 14432
rect 59284 14372 60326 14428
rect 60382 14372 60484 14428
rect 60540 14372 62528 14428
rect 62584 14372 62608 14428
rect 62664 14372 64740 14428
rect 59284 14368 64740 14372
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14428 75028 14432
rect 71284 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 75028 14428
rect 71284 14368 75028 14372
rect 964 14352 75028 14368
rect 964 14348 4740 14352
rect 964 14292 2044 14348
rect 2100 14292 4740 14348
rect 964 14288 4740 14292
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14348 10740 14352
rect 5284 14292 5540 14348
rect 5596 14292 8430 14348
rect 8486 14292 10740 14348
rect 5284 14288 10740 14292
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14348 16740 14352
rect 11284 14292 11320 14348
rect 11376 14292 14210 14348
rect 14266 14292 16740 14348
rect 11284 14288 16740 14292
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14348 17140 14352
rect 17124 14288 17140 14292
rect 17204 14288 17220 14352
rect 17284 14348 22740 14352
rect 17284 14292 19990 14348
rect 20046 14292 22740 14348
rect 17284 14288 22740 14292
rect 22804 14288 22820 14352
rect 22884 14348 22900 14352
rect 22884 14288 22900 14292
rect 22964 14288 22980 14352
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14348 28740 14352
rect 23284 14292 25770 14348
rect 25826 14292 28660 14348
rect 28716 14292 28740 14348
rect 23284 14288 28740 14292
rect 28804 14288 28820 14352
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14348 34740 14352
rect 29284 14292 31550 14348
rect 31606 14292 34440 14348
rect 34496 14292 34740 14348
rect 29284 14288 34740 14292
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14348 40740 14352
rect 35284 14292 37330 14348
rect 37386 14292 40220 14348
rect 40276 14292 40740 14348
rect 35284 14288 40740 14292
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14348 46740 14352
rect 41284 14292 43110 14348
rect 43166 14292 46000 14348
rect 46056 14292 46740 14348
rect 41284 14288 46740 14292
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14348 52740 14352
rect 47284 14292 49008 14348
rect 49064 14292 52237 14348
rect 52293 14292 52740 14348
rect 47284 14288 52740 14292
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14348 58740 14352
rect 53284 14292 53638 14348
rect 53694 14292 53806 14348
rect 53862 14292 54550 14348
rect 54606 14292 54940 14348
rect 54996 14292 55656 14348
rect 55712 14292 56234 14348
rect 56290 14292 56679 14348
rect 56735 14292 56983 14348
rect 57039 14292 57825 14348
rect 57881 14292 58465 14348
rect 58521 14292 58740 14348
rect 53284 14288 58740 14292
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14348 59060 14352
rect 59044 14292 59048 14348
rect 59044 14288 59060 14292
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14348 64740 14352
rect 59284 14292 60326 14348
rect 60382 14292 60484 14348
rect 60540 14292 62528 14348
rect 62584 14292 62608 14348
rect 62664 14292 64740 14348
rect 59284 14288 64740 14292
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14348 75028 14352
rect 71284 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 75028 14348
rect 71284 14288 75028 14292
rect 964 14264 75028 14288
rect 63718 12412 63724 12476
rect 63788 12474 63794 12476
rect 64689 12474 64755 12477
rect 63788 12472 64755 12474
rect 63788 12416 64694 12472
rect 64750 12416 64755 12472
rect 63788 12414 64755 12416
rect 63788 12412 63794 12414
rect 64689 12411 64755 12414
rect 964 12240 75028 12264
rect 964 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12236 2220 12240
rect 2284 12236 7740 12240
rect 2320 12180 5393 12236
rect 5449 12180 7740 12236
rect 2204 12176 2220 12180
rect 2284 12176 7740 12180
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12236 13740 12240
rect 8339 12180 11173 12236
rect 11229 12180 13740 12236
rect 8284 12176 13740 12180
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12176 14220 12240
rect 14284 12236 19740 12240
rect 14284 12180 16953 12236
rect 17009 12180 19740 12236
rect 14284 12176 19740 12180
rect 19804 12176 19820 12240
rect 19884 12236 19900 12240
rect 19899 12180 19900 12236
rect 19884 12176 19900 12180
rect 19964 12176 19980 12240
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12236 25740 12240
rect 20284 12180 22733 12236
rect 22789 12180 25623 12236
rect 25679 12180 25740 12236
rect 20284 12176 25740 12180
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12236 31740 12240
rect 26284 12180 28513 12236
rect 28569 12180 31403 12236
rect 31459 12180 31740 12236
rect 26284 12176 31740 12180
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12236 37740 12240
rect 32284 12180 34293 12236
rect 34349 12180 37183 12236
rect 37239 12180 37740 12236
rect 32284 12176 37740 12180
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12236 43740 12240
rect 38284 12180 40073 12236
rect 40129 12180 42963 12236
rect 43019 12180 43740 12236
rect 38284 12176 43740 12180
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12236 49740 12240
rect 44284 12180 45853 12236
rect 45909 12180 48800 12236
rect 48856 12180 49662 12236
rect 49718 12180 49740 12236
rect 44284 12176 49740 12180
rect 49804 12176 49820 12240
rect 49884 12176 49900 12240
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12236 55740 12240
rect 50284 12180 52956 12236
rect 53012 12180 53114 12236
rect 53170 12180 53470 12236
rect 53526 12180 54788 12236
rect 54844 12180 55381 12236
rect 55437 12180 55740 12236
rect 50284 12176 55740 12180
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12236 61740 12240
rect 56284 12180 56527 12236
rect 56583 12180 57963 12236
rect 58019 12180 58043 12236
rect 58099 12180 59206 12236
rect 59262 12180 59364 12236
rect 59420 12180 59672 12236
rect 59728 12180 59818 12236
rect 59874 12180 59954 12236
rect 60010 12180 60034 12236
rect 60090 12180 61740 12236
rect 56284 12176 61740 12180
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12236 67740 12240
rect 62284 12180 62326 12236
rect 62382 12180 62406 12236
rect 62462 12180 67740 12236
rect 62284 12176 67740 12180
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12236 73740 12240
rect 68284 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 73740 12236
rect 68284 12176 73740 12180
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 75028 12240
rect 964 12160 75028 12176
rect 964 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12156 2220 12160
rect 2284 12156 7740 12160
rect 2320 12100 5393 12156
rect 5449 12100 7740 12156
rect 2204 12096 2220 12100
rect 2284 12096 7740 12100
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12156 13740 12160
rect 8339 12100 11173 12156
rect 11229 12100 13740 12156
rect 8284 12096 13740 12100
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12096 14220 12160
rect 14284 12156 19740 12160
rect 14284 12100 16953 12156
rect 17009 12100 19740 12156
rect 14284 12096 19740 12100
rect 19804 12096 19820 12160
rect 19884 12156 19900 12160
rect 19899 12100 19900 12156
rect 19884 12096 19900 12100
rect 19964 12096 19980 12160
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12156 25740 12160
rect 20284 12100 22733 12156
rect 22789 12100 25623 12156
rect 25679 12100 25740 12156
rect 20284 12096 25740 12100
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12156 31740 12160
rect 26284 12100 28513 12156
rect 28569 12100 31403 12156
rect 31459 12100 31740 12156
rect 26284 12096 31740 12100
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12156 37740 12160
rect 32284 12100 34293 12156
rect 34349 12100 37183 12156
rect 37239 12100 37740 12156
rect 32284 12096 37740 12100
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12156 43740 12160
rect 38284 12100 40073 12156
rect 40129 12100 42963 12156
rect 43019 12100 43740 12156
rect 38284 12096 43740 12100
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12156 49740 12160
rect 44284 12100 45853 12156
rect 45909 12100 48800 12156
rect 48856 12100 49662 12156
rect 49718 12100 49740 12156
rect 44284 12096 49740 12100
rect 49804 12096 49820 12160
rect 49884 12096 49900 12160
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12156 55740 12160
rect 50284 12100 52956 12156
rect 53012 12100 53114 12156
rect 53170 12100 53470 12156
rect 53526 12100 54788 12156
rect 54844 12100 55381 12156
rect 55437 12100 55740 12156
rect 50284 12096 55740 12100
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12156 61740 12160
rect 56284 12100 56527 12156
rect 56583 12100 57963 12156
rect 58019 12100 58043 12156
rect 58099 12100 59206 12156
rect 59262 12100 59364 12156
rect 59420 12100 59672 12156
rect 59728 12100 59818 12156
rect 59874 12100 59954 12156
rect 60010 12100 60034 12156
rect 60090 12100 61740 12156
rect 56284 12096 61740 12100
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12156 67740 12160
rect 62284 12100 62326 12156
rect 62382 12100 62406 12156
rect 62462 12100 67740 12156
rect 62284 12096 67740 12100
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12156 73740 12160
rect 68284 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 73740 12156
rect 68284 12096 73740 12100
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 75028 12160
rect 964 12080 75028 12096
rect 964 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12076 2220 12080
rect 2284 12076 7740 12080
rect 2320 12020 5393 12076
rect 5449 12020 7740 12076
rect 2204 12016 2220 12020
rect 2284 12016 7740 12020
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12076 13740 12080
rect 8339 12020 11173 12076
rect 11229 12020 13740 12076
rect 8284 12016 13740 12020
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12016 14220 12080
rect 14284 12076 19740 12080
rect 14284 12020 16953 12076
rect 17009 12020 19740 12076
rect 14284 12016 19740 12020
rect 19804 12016 19820 12080
rect 19884 12076 19900 12080
rect 19899 12020 19900 12076
rect 19884 12016 19900 12020
rect 19964 12016 19980 12080
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12076 25740 12080
rect 20284 12020 22733 12076
rect 22789 12020 25623 12076
rect 25679 12020 25740 12076
rect 20284 12016 25740 12020
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12076 31740 12080
rect 26284 12020 28513 12076
rect 28569 12020 31403 12076
rect 31459 12020 31740 12076
rect 26284 12016 31740 12020
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12076 37740 12080
rect 32284 12020 34293 12076
rect 34349 12020 37183 12076
rect 37239 12020 37740 12076
rect 32284 12016 37740 12020
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12076 43740 12080
rect 38284 12020 40073 12076
rect 40129 12020 42963 12076
rect 43019 12020 43740 12076
rect 38284 12016 43740 12020
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12076 49740 12080
rect 44284 12020 45853 12076
rect 45909 12020 48800 12076
rect 48856 12020 49662 12076
rect 49718 12020 49740 12076
rect 44284 12016 49740 12020
rect 49804 12016 49820 12080
rect 49884 12016 49900 12080
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12076 55740 12080
rect 50284 12020 52956 12076
rect 53012 12020 53114 12076
rect 53170 12020 53470 12076
rect 53526 12020 54788 12076
rect 54844 12020 55381 12076
rect 55437 12020 55740 12076
rect 50284 12016 55740 12020
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12076 61740 12080
rect 56284 12020 56527 12076
rect 56583 12020 57963 12076
rect 58019 12020 58043 12076
rect 58099 12020 59206 12076
rect 59262 12020 59364 12076
rect 59420 12020 59672 12076
rect 59728 12020 59818 12076
rect 59874 12020 59954 12076
rect 60010 12020 60034 12076
rect 60090 12020 61740 12076
rect 56284 12016 61740 12020
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12076 67740 12080
rect 62284 12020 62326 12076
rect 62382 12020 62406 12076
rect 62462 12020 67740 12076
rect 62284 12016 67740 12020
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12076 73740 12080
rect 68284 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 73740 12076
rect 68284 12016 73740 12020
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 75028 12080
rect 964 12000 75028 12016
rect 964 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11996 2220 12000
rect 2284 11996 7740 12000
rect 2320 11940 5393 11996
rect 5449 11940 7740 11996
rect 2204 11936 2220 11940
rect 2284 11936 7740 11940
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11996 13740 12000
rect 8339 11940 11173 11996
rect 11229 11940 13740 11996
rect 8284 11936 13740 11940
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11936 14220 12000
rect 14284 11996 19740 12000
rect 14284 11940 16953 11996
rect 17009 11940 19740 11996
rect 14284 11936 19740 11940
rect 19804 11936 19820 12000
rect 19884 11996 19900 12000
rect 19899 11940 19900 11996
rect 19884 11936 19900 11940
rect 19964 11936 19980 12000
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11996 25740 12000
rect 20284 11940 22733 11996
rect 22789 11940 25623 11996
rect 25679 11940 25740 11996
rect 20284 11936 25740 11940
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11996 31740 12000
rect 26284 11940 28513 11996
rect 28569 11940 31403 11996
rect 31459 11940 31740 11996
rect 26284 11936 31740 11940
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11996 37740 12000
rect 32284 11940 34293 11996
rect 34349 11940 37183 11996
rect 37239 11940 37740 11996
rect 32284 11936 37740 11940
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11996 43740 12000
rect 38284 11940 40073 11996
rect 40129 11940 42963 11996
rect 43019 11940 43740 11996
rect 38284 11936 43740 11940
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11996 49740 12000
rect 44284 11940 45853 11996
rect 45909 11940 48800 11996
rect 48856 11940 49662 11996
rect 49718 11940 49740 11996
rect 44284 11936 49740 11940
rect 49804 11936 49820 12000
rect 49884 11936 49900 12000
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11996 55740 12000
rect 50284 11940 52956 11996
rect 53012 11940 53114 11996
rect 53170 11940 53470 11996
rect 53526 11940 54788 11996
rect 54844 11940 55381 11996
rect 55437 11940 55740 11996
rect 50284 11936 55740 11940
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11996 61740 12000
rect 56284 11940 56527 11996
rect 56583 11940 57963 11996
rect 58019 11940 58043 11996
rect 58099 11940 59206 11996
rect 59262 11940 59364 11996
rect 59420 11940 59672 11996
rect 59728 11940 59818 11996
rect 59874 11940 59954 11996
rect 60010 11940 60034 11996
rect 60090 11940 61740 11996
rect 56284 11936 61740 11940
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11996 67740 12000
rect 62284 11940 62326 11996
rect 62382 11940 62406 11996
rect 62462 11940 67740 11996
rect 62284 11936 67740 11940
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11996 73740 12000
rect 68284 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 73740 11996
rect 68284 11936 73740 11940
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 75028 12000
rect 964 11912 75028 11936
rect 63677 11796 63743 11797
rect 63677 11794 63724 11796
rect 63632 11792 63724 11794
rect 63632 11736 63682 11792
rect 63632 11734 63724 11736
rect 63677 11732 63724 11734
rect 63788 11732 63794 11796
rect 63677 11731 63743 11732
rect 65558 11596 65564 11660
rect 65628 11658 65634 11660
rect 66110 11658 66116 11660
rect 65628 11598 66116 11658
rect 65628 11596 65634 11598
rect 66110 11596 66116 11598
rect 66180 11596 66186 11660
rect 65425 11522 65491 11525
rect 65558 11522 65564 11524
rect 65425 11520 65564 11522
rect 65425 11464 65430 11520
rect 65486 11464 65564 11520
rect 65425 11462 65564 11464
rect 65425 11459 65491 11462
rect 65558 11460 65564 11462
rect 65628 11460 65634 11524
rect 30833 7714 30899 7717
rect 63902 7714 63908 7716
rect 30833 7712 63908 7714
rect 30833 7656 30838 7712
rect 30894 7656 63908 7712
rect 30833 7654 63908 7656
rect 30833 7651 30899 7654
rect 63902 7652 63908 7654
rect 63972 7652 63978 7716
rect 64965 7714 65031 7717
rect 65558 7714 65564 7716
rect 64965 7712 65564 7714
rect 64965 7656 64970 7712
rect 65026 7656 65564 7712
rect 64965 7654 65564 7656
rect 64965 7651 65031 7654
rect 65558 7652 65564 7654
rect 65628 7652 65634 7716
rect 30281 7578 30347 7581
rect 65742 7578 65748 7580
rect 30281 7576 65748 7578
rect 30281 7520 30286 7576
rect 30342 7520 65748 7576
rect 30281 7518 65748 7520
rect 30281 7515 30347 7518
rect 65742 7516 65748 7518
rect 65812 7516 65818 7580
rect 61561 7034 61627 7037
rect 61561 7032 63234 7034
rect 61561 6976 61566 7032
rect 61622 6976 63234 7032
rect 61561 6974 63234 6976
rect 61561 6971 61627 6974
rect 41045 6898 41111 6901
rect 62941 6900 63007 6901
rect 41045 6896 62682 6898
rect 41045 6840 41050 6896
rect 41106 6840 62682 6896
rect 41045 6838 62682 6840
rect 41045 6835 41111 6838
rect 29085 6762 29151 6765
rect 62622 6762 62682 6838
rect 62941 6896 62988 6900
rect 63052 6898 63058 6900
rect 63174 6898 63234 6974
rect 66662 6898 66668 6900
rect 62941 6840 62946 6896
rect 62941 6836 62988 6840
rect 63052 6838 63098 6898
rect 63174 6838 66668 6898
rect 63052 6836 63058 6838
rect 66662 6836 66668 6838
rect 66732 6836 66738 6900
rect 62941 6835 63007 6836
rect 64454 6762 64460 6764
rect 29085 6760 62498 6762
rect 29085 6704 29090 6760
rect 29146 6704 62498 6760
rect 29085 6702 62498 6704
rect 62622 6702 64460 6762
rect 29085 6699 29151 6702
rect 29729 6626 29795 6629
rect 62297 6626 62363 6629
rect 29729 6624 62363 6626
rect 29729 6568 29734 6624
rect 29790 6568 62302 6624
rect 62358 6568 62363 6624
rect 29729 6566 62363 6568
rect 62438 6626 62498 6702
rect 64454 6700 64460 6702
rect 64524 6700 64530 6764
rect 65701 6626 65767 6629
rect 62438 6624 65767 6626
rect 62438 6568 65706 6624
rect 65762 6568 65767 6624
rect 62438 6566 65767 6568
rect 29729 6563 29795 6566
rect 62297 6563 62363 6566
rect 65701 6563 65767 6566
rect 28441 6490 28507 6493
rect 65241 6490 65307 6493
rect 28441 6488 65307 6490
rect 28441 6432 28446 6488
rect 28502 6432 65246 6488
rect 65302 6432 65307 6488
rect 28441 6430 65307 6432
rect 28441 6427 28507 6430
rect 65241 6427 65307 6430
rect 55857 6354 55923 6357
rect 63953 6354 64019 6357
rect 55857 6352 64019 6354
rect 55857 6296 55862 6352
rect 55918 6296 63958 6352
rect 64014 6296 64019 6352
rect 55857 6294 64019 6296
rect 55857 6291 55923 6294
rect 63953 6291 64019 6294
rect 46749 6218 46815 6221
rect 61745 6218 61811 6221
rect 46749 6216 61811 6218
rect 46749 6160 46754 6216
rect 46810 6160 61750 6216
rect 61806 6160 61811 6216
rect 46749 6158 61811 6160
rect 46749 6155 46815 6158
rect 61745 6155 61811 6158
rect 62297 6218 62363 6221
rect 65926 6218 65932 6220
rect 62297 6216 65932 6218
rect 62297 6160 62302 6216
rect 62358 6160 65932 6216
rect 62297 6158 65932 6160
rect 62297 6155 62363 6158
rect 65926 6156 65932 6158
rect 65996 6156 66002 6220
rect 44633 6082 44699 6085
rect 55857 6082 55923 6085
rect 44633 6080 55923 6082
rect 44633 6024 44638 6080
rect 44694 6024 55862 6080
rect 55918 6024 55923 6080
rect 44633 6022 55923 6024
rect 44633 6019 44699 6022
rect 55857 6019 55923 6022
rect 59721 6082 59787 6085
rect 70393 6082 70459 6085
rect 59721 6080 70459 6082
rect 59721 6024 59726 6080
rect 59782 6024 70398 6080
rect 70454 6024 70459 6080
rect 59721 6022 70459 6024
rect 59721 6019 59787 6022
rect 70393 6019 70459 6022
rect 24577 5946 24643 5949
rect 58157 5946 58223 5949
rect 62757 5946 62823 5949
rect 24577 5944 41430 5946
rect 24577 5888 24582 5944
rect 24638 5888 41430 5944
rect 24577 5886 41430 5888
rect 24577 5883 24643 5886
rect 39982 5748 39988 5812
rect 40052 5810 40058 5812
rect 40401 5810 40467 5813
rect 40052 5808 40467 5810
rect 40052 5752 40406 5808
rect 40462 5752 40467 5808
rect 40052 5750 40467 5752
rect 41370 5810 41430 5886
rect 58157 5944 62823 5946
rect 58157 5888 58162 5944
rect 58218 5888 62762 5944
rect 62818 5888 62823 5944
rect 58157 5886 62823 5888
rect 58157 5883 58223 5886
rect 62757 5883 62823 5886
rect 61561 5810 61627 5813
rect 41370 5808 61627 5810
rect 41370 5752 61566 5808
rect 61622 5752 61627 5808
rect 41370 5750 61627 5752
rect 40052 5748 40058 5750
rect 40401 5747 40467 5750
rect 61561 5747 61627 5750
rect 61745 5810 61811 5813
rect 65977 5810 66043 5813
rect 61745 5808 66043 5810
rect 61745 5752 61750 5808
rect 61806 5752 65982 5808
rect 66038 5752 66043 5808
rect 61745 5750 66043 5752
rect 61745 5747 61811 5750
rect 65977 5747 66043 5750
rect 36997 5674 37063 5677
rect 41689 5674 41755 5677
rect 68502 5674 68508 5676
rect 36997 5672 68508 5674
rect 36997 5616 37002 5672
rect 37058 5616 41694 5672
rect 41750 5616 68508 5672
rect 36997 5614 68508 5616
rect 36997 5611 37063 5614
rect 41689 5611 41755 5614
rect 68502 5612 68508 5614
rect 68572 5612 68578 5676
rect 48957 5538 49023 5541
rect 55949 5538 56015 5541
rect 48957 5536 56015 5538
rect 48957 5480 48962 5536
rect 49018 5480 55954 5536
rect 56010 5480 56015 5536
rect 48957 5478 56015 5480
rect 48957 5475 49023 5478
rect 55949 5475 56015 5478
rect 61009 5538 61075 5541
rect 63401 5538 63467 5541
rect 61009 5536 63467 5538
rect 61009 5480 61014 5536
rect 61070 5480 63406 5536
rect 63462 5480 63467 5536
rect 61009 5478 63467 5480
rect 61009 5475 61075 5478
rect 63401 5475 63467 5478
rect 46197 5402 46263 5405
rect 64086 5402 64092 5404
rect 46197 5400 64092 5402
rect 46197 5344 46202 5400
rect 46258 5344 64092 5400
rect 46197 5342 64092 5344
rect 46197 5339 46263 5342
rect 64086 5340 64092 5342
rect 64156 5340 64162 5404
rect 27153 5266 27219 5269
rect 63309 5266 63375 5269
rect 27153 5264 63375 5266
rect 27153 5208 27158 5264
rect 27214 5208 63314 5264
rect 63370 5208 63375 5264
rect 27153 5206 63375 5208
rect 27153 5203 27219 5206
rect 63309 5203 63375 5206
rect 63585 5266 63651 5269
rect 66478 5266 66484 5268
rect 63585 5264 66484 5266
rect 63585 5208 63590 5264
rect 63646 5208 66484 5264
rect 63585 5206 66484 5208
rect 63585 5203 63651 5206
rect 66478 5204 66484 5206
rect 66548 5204 66554 5268
rect 25773 5130 25839 5133
rect 28073 5130 28139 5133
rect 25773 5128 28139 5130
rect 25773 5072 25778 5128
rect 25834 5072 28078 5128
rect 28134 5072 28139 5128
rect 25773 5070 28139 5072
rect 25773 5067 25839 5070
rect 28073 5067 28139 5070
rect 42701 5130 42767 5133
rect 64873 5130 64939 5133
rect 42701 5128 64939 5130
rect 42701 5072 42706 5128
rect 42762 5072 64878 5128
rect 64934 5072 64939 5128
rect 42701 5070 64939 5072
rect 42701 5067 42767 5070
rect 64873 5067 64939 5070
rect 27797 4994 27863 4997
rect 29729 4994 29795 4997
rect 27797 4992 29795 4994
rect 27797 4936 27802 4992
rect 27858 4936 29734 4992
rect 29790 4936 29795 4992
rect 27797 4934 29795 4936
rect 27797 4931 27863 4934
rect 29729 4931 29795 4934
rect 44725 4994 44791 4997
rect 64270 4994 64276 4996
rect 44725 4992 64276 4994
rect 44725 4936 44730 4992
rect 44786 4936 64276 4992
rect 44725 4934 64276 4936
rect 44725 4931 44791 4934
rect 64270 4932 64276 4934
rect 64340 4932 64346 4996
rect 34053 4858 34119 4861
rect 63166 4858 63172 4860
rect 34053 4856 63172 4858
rect 34053 4800 34058 4856
rect 34114 4800 63172 4856
rect 34053 4798 63172 4800
rect 34053 4795 34119 4798
rect 63166 4796 63172 4798
rect 63236 4796 63242 4860
rect 964 4592 75028 4616
rect 964 4588 4740 4592
rect 964 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4740 4588
rect 964 4528 4740 4532
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4588 16740 4592
rect 11284 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 16740 4588
rect 11284 4528 16740 4532
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4588 28740 4592
rect 23284 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 28740 4588
rect 23284 4528 28740 4532
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4588 34740 4592
rect 29284 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34740 4588
rect 29284 4528 34740 4532
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4588 46740 4592
rect 41284 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 46740 4588
rect 41284 4528 46740 4532
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4588 58740 4592
rect 53284 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 58740 4588
rect 53284 4528 58740 4532
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4588 64740 4592
rect 59284 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64740 4588
rect 59284 4528 64740 4532
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4588 75028 4592
rect 71284 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 75028 4588
rect 71284 4528 75028 4532
rect 964 4512 75028 4528
rect 964 4508 4740 4512
rect 964 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4740 4508
rect 964 4448 4740 4452
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4508 16740 4512
rect 11284 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 16740 4508
rect 11284 4448 16740 4452
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4508 28740 4512
rect 23284 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 28740 4508
rect 23284 4448 28740 4452
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4508 34740 4512
rect 29284 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34740 4508
rect 29284 4448 34740 4452
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4508 46740 4512
rect 41284 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 46740 4508
rect 41284 4448 46740 4452
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4508 58740 4512
rect 53284 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 58740 4508
rect 53284 4448 58740 4452
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4508 64740 4512
rect 59284 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64740 4508
rect 59284 4448 64740 4452
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4508 75028 4512
rect 71284 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 75028 4508
rect 71284 4448 75028 4452
rect 964 4432 75028 4448
rect 964 4428 4740 4432
rect 964 4372 4216 4428
rect 4272 4372 4296 4428
rect 4352 4372 4376 4428
rect 4432 4372 4456 4428
rect 4512 4372 4740 4428
rect 964 4368 4740 4372
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4428 16740 4432
rect 11284 4372 14216 4428
rect 14272 4372 14296 4428
rect 14352 4372 14376 4428
rect 14432 4372 14456 4428
rect 14512 4372 16740 4428
rect 11284 4368 16740 4372
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4428 28740 4432
rect 23284 4372 24216 4428
rect 24272 4372 24296 4428
rect 24352 4372 24376 4428
rect 24432 4372 24456 4428
rect 24512 4372 28740 4428
rect 23284 4368 28740 4372
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4428 34740 4432
rect 29284 4372 34216 4428
rect 34272 4372 34296 4428
rect 34352 4372 34376 4428
rect 34432 4372 34456 4428
rect 34512 4372 34740 4428
rect 29284 4368 34740 4372
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4428 46740 4432
rect 41284 4372 44216 4428
rect 44272 4372 44296 4428
rect 44352 4372 44376 4428
rect 44432 4372 44456 4428
rect 44512 4372 46740 4428
rect 41284 4368 46740 4372
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4428 58740 4432
rect 53284 4372 54216 4428
rect 54272 4372 54296 4428
rect 54352 4372 54376 4428
rect 54432 4372 54456 4428
rect 54512 4372 58740 4428
rect 53284 4368 58740 4372
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4428 64740 4432
rect 59284 4372 64216 4428
rect 64272 4372 64296 4428
rect 64352 4372 64376 4428
rect 64432 4372 64456 4428
rect 64512 4372 64740 4428
rect 59284 4368 64740 4372
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4428 75028 4432
rect 71284 4372 74216 4428
rect 74272 4372 74296 4428
rect 74352 4372 74376 4428
rect 74432 4372 74456 4428
rect 74512 4372 75028 4428
rect 71284 4368 75028 4372
rect 964 4352 75028 4368
rect 964 4348 4740 4352
rect 964 4292 4216 4348
rect 4272 4292 4296 4348
rect 4352 4292 4376 4348
rect 4432 4292 4456 4348
rect 4512 4292 4740 4348
rect 964 4288 4740 4292
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4348 16740 4352
rect 11284 4292 14216 4348
rect 14272 4292 14296 4348
rect 14352 4292 14376 4348
rect 14432 4292 14456 4348
rect 14512 4292 16740 4348
rect 11284 4288 16740 4292
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4348 28740 4352
rect 23284 4292 24216 4348
rect 24272 4292 24296 4348
rect 24352 4292 24376 4348
rect 24432 4292 24456 4348
rect 24512 4292 28740 4348
rect 23284 4288 28740 4292
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4348 34740 4352
rect 29284 4292 34216 4348
rect 34272 4292 34296 4348
rect 34352 4292 34376 4348
rect 34432 4292 34456 4348
rect 34512 4292 34740 4348
rect 29284 4288 34740 4292
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4348 46740 4352
rect 41284 4292 44216 4348
rect 44272 4292 44296 4348
rect 44352 4292 44376 4348
rect 44432 4292 44456 4348
rect 44512 4292 46740 4348
rect 41284 4288 46740 4292
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4348 58740 4352
rect 53284 4292 54216 4348
rect 54272 4292 54296 4348
rect 54352 4292 54376 4348
rect 54432 4292 54456 4348
rect 54512 4292 58740 4348
rect 53284 4288 58740 4292
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4348 64740 4352
rect 59284 4292 64216 4348
rect 64272 4292 64296 4348
rect 64352 4292 64376 4348
rect 64432 4292 64456 4348
rect 64512 4292 64740 4348
rect 59284 4288 64740 4292
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4348 75028 4352
rect 71284 4292 74216 4348
rect 74272 4292 74296 4348
rect 74352 4292 74376 4348
rect 74432 4292 74456 4348
rect 74512 4292 75028 4348
rect 71284 4288 75028 4292
rect 964 4264 75028 4288
rect 43345 4178 43411 4181
rect 44725 4178 44791 4181
rect 43345 4176 44791 4178
rect 43345 4120 43350 4176
rect 43406 4120 44730 4176
rect 44786 4120 44791 4176
rect 43345 4118 44791 4120
rect 43345 4115 43411 4118
rect 44725 4115 44791 4118
rect 60641 4178 60707 4181
rect 61377 4178 61443 4181
rect 60641 4176 61443 4178
rect 60641 4120 60646 4176
rect 60702 4120 61382 4176
rect 61438 4120 61443 4176
rect 60641 4118 61443 4120
rect 60641 4115 60707 4118
rect 61377 4115 61443 4118
rect 31293 4042 31359 4045
rect 66110 4042 66116 4044
rect 31293 4040 66116 4042
rect 31293 3984 31298 4040
rect 31354 3984 66116 4040
rect 31293 3982 66116 3984
rect 31293 3979 31359 3982
rect 66110 3980 66116 3982
rect 66180 3980 66186 4044
rect 14733 3362 14799 3365
rect 39982 3362 39988 3364
rect 14733 3360 39988 3362
rect 14733 3304 14738 3360
rect 14794 3304 39988 3360
rect 14733 3302 39988 3304
rect 14733 3299 14799 3302
rect 39982 3300 39988 3302
rect 40052 3300 40058 3364
rect 41413 3362 41479 3365
rect 66294 3362 66300 3364
rect 41413 3360 66300 3362
rect 41413 3304 41418 3360
rect 41474 3304 66300 3360
rect 41413 3302 66300 3304
rect 41413 3299 41479 3302
rect 66294 3300 66300 3302
rect 66364 3300 66370 3364
rect 20897 3226 20963 3229
rect 25865 3226 25931 3229
rect 20897 3224 25931 3226
rect 20897 3168 20902 3224
rect 20958 3168 25870 3224
rect 25926 3168 25931 3224
rect 20897 3166 25931 3168
rect 20897 3163 20963 3166
rect 25865 3163 25931 3166
rect 26141 3090 26207 3093
rect 28901 3090 28967 3093
rect 26141 3088 28967 3090
rect 26141 3032 26146 3088
rect 26202 3032 28906 3088
rect 28962 3032 28967 3088
rect 26141 3030 28967 3032
rect 26141 3027 26207 3030
rect 28901 3027 28967 3030
rect 32213 3090 32279 3093
rect 63585 3090 63651 3093
rect 32213 3088 63651 3090
rect 32213 3032 32218 3088
rect 32274 3032 63590 3088
rect 63646 3032 63651 3088
rect 32213 3030 63651 3032
rect 32213 3027 32279 3030
rect 63585 3027 63651 3030
rect 964 2240 75028 2264
rect 964 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2236 1900 2240
rect 1964 2236 1980 2240
rect 2044 2236 2060 2240
rect 2124 2236 2140 2240
rect 1884 2176 1900 2180
rect 1964 2176 1980 2180
rect 2044 2176 2060 2180
rect 2124 2176 2140 2180
rect 2204 2176 2220 2240
rect 2284 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2236 13740 2240
rect 8284 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 13740 2236
rect 8284 2176 13740 2180
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2236 25740 2240
rect 20284 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 25740 2236
rect 20284 2176 25740 2180
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2236 31900 2240
rect 31964 2236 31980 2240
rect 32044 2236 32060 2240
rect 32124 2236 32140 2240
rect 31884 2176 31900 2180
rect 31964 2176 31980 2180
rect 32044 2176 32060 2180
rect 32124 2176 32140 2180
rect 32204 2176 32220 2240
rect 32284 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2236 43740 2240
rect 38284 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 43740 2236
rect 38284 2176 43740 2180
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2236 55740 2240
rect 50284 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 55740 2236
rect 50284 2176 55740 2180
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2236 61900 2240
rect 61964 2236 61980 2240
rect 62044 2236 62060 2240
rect 62124 2236 62140 2240
rect 61884 2176 61900 2180
rect 61964 2176 61980 2180
rect 62044 2176 62060 2180
rect 62124 2176 62140 2180
rect 62204 2176 62220 2240
rect 62284 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2236 73740 2240
rect 68284 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 73740 2236
rect 68284 2176 73740 2180
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 75028 2240
rect 964 2160 75028 2176
rect 964 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2156 1900 2160
rect 1964 2156 1980 2160
rect 2044 2156 2060 2160
rect 2124 2156 2140 2160
rect 1884 2096 1900 2100
rect 1964 2096 1980 2100
rect 2044 2096 2060 2100
rect 2124 2096 2140 2100
rect 2204 2096 2220 2160
rect 2284 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2156 13740 2160
rect 8284 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 13740 2156
rect 8284 2096 13740 2100
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2156 25740 2160
rect 20284 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 25740 2156
rect 20284 2096 25740 2100
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2156 31900 2160
rect 31964 2156 31980 2160
rect 32044 2156 32060 2160
rect 32124 2156 32140 2160
rect 31884 2096 31900 2100
rect 31964 2096 31980 2100
rect 32044 2096 32060 2100
rect 32124 2096 32140 2100
rect 32204 2096 32220 2160
rect 32284 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2156 43740 2160
rect 38284 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 43740 2156
rect 38284 2096 43740 2100
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2156 55740 2160
rect 50284 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 55740 2156
rect 50284 2096 55740 2100
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2156 61900 2160
rect 61964 2156 61980 2160
rect 62044 2156 62060 2160
rect 62124 2156 62140 2160
rect 61884 2096 61900 2100
rect 61964 2096 61980 2100
rect 62044 2096 62060 2100
rect 62124 2096 62140 2100
rect 62204 2096 62220 2160
rect 62284 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2156 73740 2160
rect 68284 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 73740 2156
rect 68284 2096 73740 2100
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 75028 2160
rect 964 2080 75028 2096
rect 964 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2076 1900 2080
rect 1964 2076 1980 2080
rect 2044 2076 2060 2080
rect 2124 2076 2140 2080
rect 1884 2016 1900 2020
rect 1964 2016 1980 2020
rect 2044 2016 2060 2020
rect 2124 2016 2140 2020
rect 2204 2016 2220 2080
rect 2284 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2076 13740 2080
rect 8284 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 13740 2076
rect 8284 2016 13740 2020
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2076 25740 2080
rect 20284 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 25740 2076
rect 20284 2016 25740 2020
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2076 31900 2080
rect 31964 2076 31980 2080
rect 32044 2076 32060 2080
rect 32124 2076 32140 2080
rect 31884 2016 31900 2020
rect 31964 2016 31980 2020
rect 32044 2016 32060 2020
rect 32124 2016 32140 2020
rect 32204 2016 32220 2080
rect 32284 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2076 43740 2080
rect 38284 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 43740 2076
rect 38284 2016 43740 2020
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2076 55740 2080
rect 50284 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 55740 2076
rect 50284 2016 55740 2020
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2076 61900 2080
rect 61964 2076 61980 2080
rect 62044 2076 62060 2080
rect 62124 2076 62140 2080
rect 61884 2016 61900 2020
rect 61964 2016 61980 2020
rect 62044 2016 62060 2020
rect 62124 2016 62140 2020
rect 62204 2016 62220 2080
rect 62284 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2076 73740 2080
rect 68284 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 73740 2076
rect 68284 2016 73740 2020
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 75028 2080
rect 964 2000 75028 2016
rect 964 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1996 1900 2000
rect 1964 1996 1980 2000
rect 2044 1996 2060 2000
rect 2124 1996 2140 2000
rect 1884 1936 1900 1940
rect 1964 1936 1980 1940
rect 2044 1936 2060 1940
rect 2124 1936 2140 1940
rect 2204 1936 2220 2000
rect 2284 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1996 13740 2000
rect 8284 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 13740 1996
rect 8284 1936 13740 1940
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1996 25740 2000
rect 20284 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 25740 1996
rect 20284 1936 25740 1940
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1996 31900 2000
rect 31964 1996 31980 2000
rect 32044 1996 32060 2000
rect 32124 1996 32140 2000
rect 31884 1936 31900 1940
rect 31964 1936 31980 1940
rect 32044 1936 32060 1940
rect 32124 1936 32140 1940
rect 32204 1936 32220 2000
rect 32284 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1996 43740 2000
rect 38284 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 43740 1996
rect 38284 1936 43740 1940
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1996 55740 2000
rect 50284 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 55740 1996
rect 50284 1936 55740 1940
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1996 61900 2000
rect 61964 1996 61980 2000
rect 62044 1996 62060 2000
rect 62124 1996 62140 2000
rect 61884 1936 61900 1940
rect 61964 1936 61980 1940
rect 62044 1936 62060 1940
rect 62124 1936 62140 1940
rect 62204 1936 62220 2000
rect 62284 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1996 73740 2000
rect 68284 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 73740 1996
rect 68284 1936 73740 1940
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 75028 2000
rect 964 1912 75028 1936
rect 31109 1594 31175 1597
rect 35985 1594 36051 1597
rect 31109 1592 36051 1594
rect 31109 1536 31114 1592
rect 31170 1536 35990 1592
rect 36046 1536 36051 1592
rect 31109 1534 36051 1536
rect 31109 1531 31175 1534
rect 35985 1531 36051 1534
rect 23197 1458 23263 1461
rect 28441 1458 28507 1461
rect 23197 1456 28507 1458
rect 23197 1400 23202 1456
rect 23258 1400 28446 1456
rect 28502 1400 28507 1456
rect 23197 1398 28507 1400
rect 23197 1395 23263 1398
rect 28441 1395 28507 1398
<< via3 >>
rect 4740 84528 4804 84592
rect 4820 84528 4884 84592
rect 4900 84528 4964 84592
rect 4980 84528 5044 84592
rect 5060 84528 5124 84592
rect 5140 84528 5204 84592
rect 5220 84528 5284 84592
rect 10740 84528 10804 84592
rect 10820 84528 10884 84592
rect 10900 84528 10964 84592
rect 10980 84528 11044 84592
rect 11060 84528 11124 84592
rect 11140 84528 11204 84592
rect 11220 84528 11284 84592
rect 16740 84528 16804 84592
rect 16820 84528 16884 84592
rect 16900 84528 16964 84592
rect 16980 84528 17044 84592
rect 17060 84588 17124 84592
rect 17140 84588 17204 84592
rect 17060 84532 17100 84588
rect 17100 84532 17124 84588
rect 17140 84532 17156 84588
rect 17156 84532 17204 84588
rect 17060 84528 17124 84532
rect 17140 84528 17204 84532
rect 17220 84528 17284 84592
rect 22740 84528 22804 84592
rect 22820 84588 22884 84592
rect 22900 84588 22964 84592
rect 22820 84532 22880 84588
rect 22880 84532 22884 84588
rect 22900 84532 22936 84588
rect 22936 84532 22964 84588
rect 22820 84528 22884 84532
rect 22900 84528 22964 84532
rect 22980 84528 23044 84592
rect 23060 84528 23124 84592
rect 23140 84528 23204 84592
rect 23220 84528 23284 84592
rect 28740 84528 28804 84592
rect 28820 84528 28884 84592
rect 28900 84528 28964 84592
rect 28980 84528 29044 84592
rect 29060 84528 29124 84592
rect 29140 84528 29204 84592
rect 29220 84528 29284 84592
rect 34740 84528 34804 84592
rect 34820 84528 34884 84592
rect 34900 84528 34964 84592
rect 34980 84528 35044 84592
rect 35060 84528 35124 84592
rect 35140 84528 35204 84592
rect 35220 84528 35284 84592
rect 40740 84528 40804 84592
rect 40820 84528 40884 84592
rect 40900 84528 40964 84592
rect 40980 84528 41044 84592
rect 41060 84528 41124 84592
rect 41140 84528 41204 84592
rect 41220 84528 41284 84592
rect 46740 84528 46804 84592
rect 46820 84528 46884 84592
rect 46900 84528 46964 84592
rect 46980 84528 47044 84592
rect 47060 84528 47124 84592
rect 47140 84528 47204 84592
rect 47220 84528 47284 84592
rect 52740 84528 52804 84592
rect 52820 84528 52884 84592
rect 52900 84528 52964 84592
rect 52980 84528 53044 84592
rect 53060 84528 53124 84592
rect 53140 84528 53204 84592
rect 53220 84528 53284 84592
rect 58740 84528 58804 84592
rect 58820 84528 58884 84592
rect 58900 84528 58964 84592
rect 58980 84528 59044 84592
rect 59060 84588 59124 84592
rect 59060 84532 59104 84588
rect 59104 84532 59124 84588
rect 59060 84528 59124 84532
rect 59140 84528 59204 84592
rect 59220 84528 59284 84592
rect 64740 84528 64804 84592
rect 64820 84528 64884 84592
rect 64900 84528 64964 84592
rect 64980 84528 65044 84592
rect 65060 84528 65124 84592
rect 65140 84528 65204 84592
rect 65220 84528 65284 84592
rect 70740 84528 70804 84592
rect 70820 84528 70884 84592
rect 70900 84528 70964 84592
rect 70980 84528 71044 84592
rect 71060 84528 71124 84592
rect 71140 84528 71204 84592
rect 71220 84528 71284 84592
rect 4740 84448 4804 84512
rect 4820 84448 4884 84512
rect 4900 84448 4964 84512
rect 4980 84448 5044 84512
rect 5060 84448 5124 84512
rect 5140 84448 5204 84512
rect 5220 84448 5284 84512
rect 10740 84448 10804 84512
rect 10820 84448 10884 84512
rect 10900 84448 10964 84512
rect 10980 84448 11044 84512
rect 11060 84448 11124 84512
rect 11140 84448 11204 84512
rect 11220 84448 11284 84512
rect 16740 84448 16804 84512
rect 16820 84448 16884 84512
rect 16900 84448 16964 84512
rect 16980 84448 17044 84512
rect 17060 84508 17124 84512
rect 17140 84508 17204 84512
rect 17060 84452 17100 84508
rect 17100 84452 17124 84508
rect 17140 84452 17156 84508
rect 17156 84452 17204 84508
rect 17060 84448 17124 84452
rect 17140 84448 17204 84452
rect 17220 84448 17284 84512
rect 22740 84448 22804 84512
rect 22820 84508 22884 84512
rect 22900 84508 22964 84512
rect 22820 84452 22880 84508
rect 22880 84452 22884 84508
rect 22900 84452 22936 84508
rect 22936 84452 22964 84508
rect 22820 84448 22884 84452
rect 22900 84448 22964 84452
rect 22980 84448 23044 84512
rect 23060 84448 23124 84512
rect 23140 84448 23204 84512
rect 23220 84448 23284 84512
rect 28740 84448 28804 84512
rect 28820 84448 28884 84512
rect 28900 84448 28964 84512
rect 28980 84448 29044 84512
rect 29060 84448 29124 84512
rect 29140 84448 29204 84512
rect 29220 84448 29284 84512
rect 34740 84448 34804 84512
rect 34820 84448 34884 84512
rect 34900 84448 34964 84512
rect 34980 84448 35044 84512
rect 35060 84448 35124 84512
rect 35140 84448 35204 84512
rect 35220 84448 35284 84512
rect 40740 84448 40804 84512
rect 40820 84448 40884 84512
rect 40900 84448 40964 84512
rect 40980 84448 41044 84512
rect 41060 84448 41124 84512
rect 41140 84448 41204 84512
rect 41220 84448 41284 84512
rect 46740 84448 46804 84512
rect 46820 84448 46884 84512
rect 46900 84448 46964 84512
rect 46980 84448 47044 84512
rect 47060 84448 47124 84512
rect 47140 84448 47204 84512
rect 47220 84448 47284 84512
rect 52740 84448 52804 84512
rect 52820 84448 52884 84512
rect 52900 84448 52964 84512
rect 52980 84448 53044 84512
rect 53060 84448 53124 84512
rect 53140 84448 53204 84512
rect 53220 84448 53284 84512
rect 58740 84448 58804 84512
rect 58820 84448 58884 84512
rect 58900 84448 58964 84512
rect 58980 84448 59044 84512
rect 59060 84508 59124 84512
rect 59060 84452 59104 84508
rect 59104 84452 59124 84508
rect 59060 84448 59124 84452
rect 59140 84448 59204 84512
rect 59220 84448 59284 84512
rect 64740 84448 64804 84512
rect 64820 84448 64884 84512
rect 64900 84448 64964 84512
rect 64980 84448 65044 84512
rect 65060 84448 65124 84512
rect 65140 84448 65204 84512
rect 65220 84448 65284 84512
rect 70740 84448 70804 84512
rect 70820 84448 70884 84512
rect 70900 84448 70964 84512
rect 70980 84448 71044 84512
rect 71060 84448 71124 84512
rect 71140 84448 71204 84512
rect 71220 84448 71284 84512
rect 4740 84368 4804 84432
rect 4820 84368 4884 84432
rect 4900 84368 4964 84432
rect 4980 84368 5044 84432
rect 5060 84368 5124 84432
rect 5140 84368 5204 84432
rect 5220 84368 5284 84432
rect 10740 84368 10804 84432
rect 10820 84368 10884 84432
rect 10900 84368 10964 84432
rect 10980 84368 11044 84432
rect 11060 84368 11124 84432
rect 11140 84368 11204 84432
rect 11220 84368 11284 84432
rect 16740 84368 16804 84432
rect 16820 84368 16884 84432
rect 16900 84368 16964 84432
rect 16980 84368 17044 84432
rect 17060 84428 17124 84432
rect 17140 84428 17204 84432
rect 17060 84372 17100 84428
rect 17100 84372 17124 84428
rect 17140 84372 17156 84428
rect 17156 84372 17204 84428
rect 17060 84368 17124 84372
rect 17140 84368 17204 84372
rect 17220 84368 17284 84432
rect 22740 84368 22804 84432
rect 22820 84428 22884 84432
rect 22900 84428 22964 84432
rect 22820 84372 22880 84428
rect 22880 84372 22884 84428
rect 22900 84372 22936 84428
rect 22936 84372 22964 84428
rect 22820 84368 22884 84372
rect 22900 84368 22964 84372
rect 22980 84368 23044 84432
rect 23060 84368 23124 84432
rect 23140 84368 23204 84432
rect 23220 84368 23284 84432
rect 28740 84368 28804 84432
rect 28820 84368 28884 84432
rect 28900 84368 28964 84432
rect 28980 84368 29044 84432
rect 29060 84368 29124 84432
rect 29140 84368 29204 84432
rect 29220 84368 29284 84432
rect 34740 84368 34804 84432
rect 34820 84368 34884 84432
rect 34900 84368 34964 84432
rect 34980 84368 35044 84432
rect 35060 84368 35124 84432
rect 35140 84368 35204 84432
rect 35220 84368 35284 84432
rect 40740 84368 40804 84432
rect 40820 84368 40884 84432
rect 40900 84368 40964 84432
rect 40980 84368 41044 84432
rect 41060 84368 41124 84432
rect 41140 84368 41204 84432
rect 41220 84368 41284 84432
rect 46740 84368 46804 84432
rect 46820 84368 46884 84432
rect 46900 84368 46964 84432
rect 46980 84368 47044 84432
rect 47060 84368 47124 84432
rect 47140 84368 47204 84432
rect 47220 84368 47284 84432
rect 52740 84368 52804 84432
rect 52820 84368 52884 84432
rect 52900 84368 52964 84432
rect 52980 84368 53044 84432
rect 53060 84368 53124 84432
rect 53140 84368 53204 84432
rect 53220 84368 53284 84432
rect 58740 84368 58804 84432
rect 58820 84368 58884 84432
rect 58900 84368 58964 84432
rect 58980 84368 59044 84432
rect 59060 84428 59124 84432
rect 59060 84372 59104 84428
rect 59104 84372 59124 84428
rect 59060 84368 59124 84372
rect 59140 84368 59204 84432
rect 59220 84368 59284 84432
rect 64740 84368 64804 84432
rect 64820 84368 64884 84432
rect 64900 84368 64964 84432
rect 64980 84368 65044 84432
rect 65060 84368 65124 84432
rect 65140 84368 65204 84432
rect 65220 84368 65284 84432
rect 70740 84368 70804 84432
rect 70820 84368 70884 84432
rect 70900 84368 70964 84432
rect 70980 84368 71044 84432
rect 71060 84368 71124 84432
rect 71140 84368 71204 84432
rect 71220 84368 71284 84432
rect 4740 84288 4804 84352
rect 4820 84288 4884 84352
rect 4900 84288 4964 84352
rect 4980 84288 5044 84352
rect 5060 84288 5124 84352
rect 5140 84288 5204 84352
rect 5220 84288 5284 84352
rect 10740 84288 10804 84352
rect 10820 84288 10884 84352
rect 10900 84288 10964 84352
rect 10980 84288 11044 84352
rect 11060 84288 11124 84352
rect 11140 84288 11204 84352
rect 11220 84288 11284 84352
rect 16740 84288 16804 84352
rect 16820 84288 16884 84352
rect 16900 84288 16964 84352
rect 16980 84288 17044 84352
rect 17060 84348 17124 84352
rect 17140 84348 17204 84352
rect 17060 84292 17100 84348
rect 17100 84292 17124 84348
rect 17140 84292 17156 84348
rect 17156 84292 17204 84348
rect 17060 84288 17124 84292
rect 17140 84288 17204 84292
rect 17220 84288 17284 84352
rect 22740 84288 22804 84352
rect 22820 84348 22884 84352
rect 22900 84348 22964 84352
rect 22820 84292 22880 84348
rect 22880 84292 22884 84348
rect 22900 84292 22936 84348
rect 22936 84292 22964 84348
rect 22820 84288 22884 84292
rect 22900 84288 22964 84292
rect 22980 84288 23044 84352
rect 23060 84288 23124 84352
rect 23140 84288 23204 84352
rect 23220 84288 23284 84352
rect 28740 84288 28804 84352
rect 28820 84288 28884 84352
rect 28900 84288 28964 84352
rect 28980 84288 29044 84352
rect 29060 84288 29124 84352
rect 29140 84288 29204 84352
rect 29220 84288 29284 84352
rect 34740 84288 34804 84352
rect 34820 84288 34884 84352
rect 34900 84288 34964 84352
rect 34980 84288 35044 84352
rect 35060 84288 35124 84352
rect 35140 84288 35204 84352
rect 35220 84288 35284 84352
rect 40740 84288 40804 84352
rect 40820 84288 40884 84352
rect 40900 84288 40964 84352
rect 40980 84288 41044 84352
rect 41060 84288 41124 84352
rect 41140 84288 41204 84352
rect 41220 84288 41284 84352
rect 46740 84288 46804 84352
rect 46820 84288 46884 84352
rect 46900 84288 46964 84352
rect 46980 84288 47044 84352
rect 47060 84288 47124 84352
rect 47140 84288 47204 84352
rect 47220 84288 47284 84352
rect 52740 84288 52804 84352
rect 52820 84288 52884 84352
rect 52900 84288 52964 84352
rect 52980 84288 53044 84352
rect 53060 84288 53124 84352
rect 53140 84288 53204 84352
rect 53220 84288 53284 84352
rect 58740 84288 58804 84352
rect 58820 84288 58884 84352
rect 58900 84288 58964 84352
rect 58980 84288 59044 84352
rect 59060 84348 59124 84352
rect 59060 84292 59104 84348
rect 59104 84292 59124 84348
rect 59060 84288 59124 84292
rect 59140 84288 59204 84352
rect 59220 84288 59284 84352
rect 64740 84288 64804 84352
rect 64820 84288 64884 84352
rect 64900 84288 64964 84352
rect 64980 84288 65044 84352
rect 65060 84288 65124 84352
rect 65140 84288 65204 84352
rect 65220 84288 65284 84352
rect 70740 84288 70804 84352
rect 70820 84288 70884 84352
rect 70900 84288 70964 84352
rect 70980 84288 71044 84352
rect 71060 84288 71124 84352
rect 71140 84288 71204 84352
rect 71220 84288 71284 84352
rect 1740 82176 1804 82240
rect 1820 82176 1884 82240
rect 1900 82176 1964 82240
rect 1980 82176 2044 82240
rect 2060 82176 2124 82240
rect 2140 82236 2204 82240
rect 2220 82236 2284 82240
rect 2140 82180 2184 82236
rect 2184 82180 2204 82236
rect 2220 82180 2240 82236
rect 2240 82180 2264 82236
rect 2264 82180 2284 82236
rect 2140 82176 2204 82180
rect 2220 82176 2284 82180
rect 7740 82176 7804 82240
rect 7820 82176 7884 82240
rect 7900 82176 7964 82240
rect 7980 82176 8044 82240
rect 8060 82176 8124 82240
rect 8140 82176 8204 82240
rect 8220 82236 8284 82240
rect 8220 82180 8283 82236
rect 8283 82180 8284 82236
rect 8220 82176 8284 82180
rect 13740 82176 13804 82240
rect 13820 82176 13884 82240
rect 13900 82176 13964 82240
rect 13980 82176 14044 82240
rect 14060 82236 14124 82240
rect 14060 82180 14063 82236
rect 14063 82180 14119 82236
rect 14119 82180 14124 82236
rect 14060 82176 14124 82180
rect 14140 82176 14204 82240
rect 14220 82176 14284 82240
rect 19740 82176 19804 82240
rect 19820 82236 19884 82240
rect 19820 82180 19843 82236
rect 19843 82180 19884 82236
rect 19820 82176 19884 82180
rect 19900 82176 19964 82240
rect 19980 82176 20044 82240
rect 20060 82176 20124 82240
rect 20140 82176 20204 82240
rect 20220 82176 20284 82240
rect 25740 82176 25804 82240
rect 25820 82176 25884 82240
rect 25900 82176 25964 82240
rect 25980 82176 26044 82240
rect 26060 82176 26124 82240
rect 26140 82176 26204 82240
rect 26220 82176 26284 82240
rect 31740 82176 31804 82240
rect 31820 82176 31884 82240
rect 31900 82176 31964 82240
rect 31980 82176 32044 82240
rect 32060 82176 32124 82240
rect 32140 82176 32204 82240
rect 32220 82176 32284 82240
rect 37740 82176 37804 82240
rect 37820 82176 37884 82240
rect 37900 82176 37964 82240
rect 37980 82176 38044 82240
rect 38060 82176 38124 82240
rect 38140 82176 38204 82240
rect 38220 82176 38284 82240
rect 43740 82176 43804 82240
rect 43820 82176 43884 82240
rect 43900 82176 43964 82240
rect 43980 82176 44044 82240
rect 44060 82176 44124 82240
rect 44140 82176 44204 82240
rect 44220 82176 44284 82240
rect 49740 82236 49804 82240
rect 49740 82180 49742 82236
rect 49742 82180 49798 82236
rect 49798 82180 49804 82236
rect 49740 82176 49804 82180
rect 49820 82176 49884 82240
rect 49900 82176 49964 82240
rect 49980 82176 50044 82240
rect 50060 82176 50124 82240
rect 50140 82176 50204 82240
rect 50220 82176 50284 82240
rect 55740 82176 55804 82240
rect 55820 82176 55884 82240
rect 55900 82176 55964 82240
rect 55980 82176 56044 82240
rect 56060 82176 56124 82240
rect 56140 82176 56204 82240
rect 56220 82176 56284 82240
rect 61740 82176 61804 82240
rect 61820 82176 61884 82240
rect 61900 82176 61964 82240
rect 61980 82176 62044 82240
rect 62060 82176 62124 82240
rect 62140 82176 62204 82240
rect 62220 82176 62284 82240
rect 67740 82176 67804 82240
rect 67820 82176 67884 82240
rect 67900 82176 67964 82240
rect 67980 82176 68044 82240
rect 68060 82176 68124 82240
rect 68140 82176 68204 82240
rect 68220 82176 68284 82240
rect 73740 82176 73804 82240
rect 73820 82176 73884 82240
rect 73900 82176 73964 82240
rect 73980 82176 74044 82240
rect 74060 82176 74124 82240
rect 74140 82176 74204 82240
rect 74220 82176 74284 82240
rect 1740 82096 1804 82160
rect 1820 82096 1884 82160
rect 1900 82096 1964 82160
rect 1980 82096 2044 82160
rect 2060 82096 2124 82160
rect 2140 82156 2204 82160
rect 2220 82156 2284 82160
rect 2140 82100 2184 82156
rect 2184 82100 2204 82156
rect 2220 82100 2240 82156
rect 2240 82100 2264 82156
rect 2264 82100 2284 82156
rect 2140 82096 2204 82100
rect 2220 82096 2284 82100
rect 7740 82096 7804 82160
rect 7820 82096 7884 82160
rect 7900 82096 7964 82160
rect 7980 82096 8044 82160
rect 8060 82096 8124 82160
rect 8140 82096 8204 82160
rect 8220 82156 8284 82160
rect 8220 82100 8283 82156
rect 8283 82100 8284 82156
rect 8220 82096 8284 82100
rect 13740 82096 13804 82160
rect 13820 82096 13884 82160
rect 13900 82096 13964 82160
rect 13980 82096 14044 82160
rect 14060 82156 14124 82160
rect 14060 82100 14063 82156
rect 14063 82100 14119 82156
rect 14119 82100 14124 82156
rect 14060 82096 14124 82100
rect 14140 82096 14204 82160
rect 14220 82096 14284 82160
rect 19740 82096 19804 82160
rect 19820 82156 19884 82160
rect 19820 82100 19843 82156
rect 19843 82100 19884 82156
rect 19820 82096 19884 82100
rect 19900 82096 19964 82160
rect 19980 82096 20044 82160
rect 20060 82096 20124 82160
rect 20140 82096 20204 82160
rect 20220 82096 20284 82160
rect 25740 82096 25804 82160
rect 25820 82096 25884 82160
rect 25900 82096 25964 82160
rect 25980 82096 26044 82160
rect 26060 82096 26124 82160
rect 26140 82096 26204 82160
rect 26220 82096 26284 82160
rect 31740 82096 31804 82160
rect 31820 82096 31884 82160
rect 31900 82096 31964 82160
rect 31980 82096 32044 82160
rect 32060 82096 32124 82160
rect 32140 82096 32204 82160
rect 32220 82096 32284 82160
rect 37740 82096 37804 82160
rect 37820 82096 37884 82160
rect 37900 82096 37964 82160
rect 37980 82096 38044 82160
rect 38060 82096 38124 82160
rect 38140 82096 38204 82160
rect 38220 82096 38284 82160
rect 43740 82096 43804 82160
rect 43820 82096 43884 82160
rect 43900 82096 43964 82160
rect 43980 82096 44044 82160
rect 44060 82096 44124 82160
rect 44140 82096 44204 82160
rect 44220 82096 44284 82160
rect 49740 82156 49804 82160
rect 49740 82100 49742 82156
rect 49742 82100 49798 82156
rect 49798 82100 49804 82156
rect 49740 82096 49804 82100
rect 49820 82096 49884 82160
rect 49900 82096 49964 82160
rect 49980 82096 50044 82160
rect 50060 82096 50124 82160
rect 50140 82096 50204 82160
rect 50220 82096 50284 82160
rect 55740 82096 55804 82160
rect 55820 82096 55884 82160
rect 55900 82096 55964 82160
rect 55980 82096 56044 82160
rect 56060 82096 56124 82160
rect 56140 82096 56204 82160
rect 56220 82096 56284 82160
rect 61740 82096 61804 82160
rect 61820 82096 61884 82160
rect 61900 82096 61964 82160
rect 61980 82096 62044 82160
rect 62060 82096 62124 82160
rect 62140 82096 62204 82160
rect 62220 82096 62284 82160
rect 67740 82096 67804 82160
rect 67820 82096 67884 82160
rect 67900 82096 67964 82160
rect 67980 82096 68044 82160
rect 68060 82096 68124 82160
rect 68140 82096 68204 82160
rect 68220 82096 68284 82160
rect 73740 82096 73804 82160
rect 73820 82096 73884 82160
rect 73900 82096 73964 82160
rect 73980 82096 74044 82160
rect 74060 82096 74124 82160
rect 74140 82096 74204 82160
rect 74220 82096 74284 82160
rect 1740 82016 1804 82080
rect 1820 82016 1884 82080
rect 1900 82016 1964 82080
rect 1980 82016 2044 82080
rect 2060 82016 2124 82080
rect 2140 82076 2204 82080
rect 2220 82076 2284 82080
rect 2140 82020 2184 82076
rect 2184 82020 2204 82076
rect 2220 82020 2240 82076
rect 2240 82020 2264 82076
rect 2264 82020 2284 82076
rect 2140 82016 2204 82020
rect 2220 82016 2284 82020
rect 7740 82016 7804 82080
rect 7820 82016 7884 82080
rect 7900 82016 7964 82080
rect 7980 82016 8044 82080
rect 8060 82016 8124 82080
rect 8140 82016 8204 82080
rect 8220 82076 8284 82080
rect 8220 82020 8283 82076
rect 8283 82020 8284 82076
rect 8220 82016 8284 82020
rect 13740 82016 13804 82080
rect 13820 82016 13884 82080
rect 13900 82016 13964 82080
rect 13980 82016 14044 82080
rect 14060 82076 14124 82080
rect 14060 82020 14063 82076
rect 14063 82020 14119 82076
rect 14119 82020 14124 82076
rect 14060 82016 14124 82020
rect 14140 82016 14204 82080
rect 14220 82016 14284 82080
rect 19740 82016 19804 82080
rect 19820 82076 19884 82080
rect 19820 82020 19843 82076
rect 19843 82020 19884 82076
rect 19820 82016 19884 82020
rect 19900 82016 19964 82080
rect 19980 82016 20044 82080
rect 20060 82016 20124 82080
rect 20140 82016 20204 82080
rect 20220 82016 20284 82080
rect 25740 82016 25804 82080
rect 25820 82016 25884 82080
rect 25900 82016 25964 82080
rect 25980 82016 26044 82080
rect 26060 82016 26124 82080
rect 26140 82016 26204 82080
rect 26220 82016 26284 82080
rect 31740 82016 31804 82080
rect 31820 82016 31884 82080
rect 31900 82016 31964 82080
rect 31980 82016 32044 82080
rect 32060 82016 32124 82080
rect 32140 82016 32204 82080
rect 32220 82016 32284 82080
rect 37740 82016 37804 82080
rect 37820 82016 37884 82080
rect 37900 82016 37964 82080
rect 37980 82016 38044 82080
rect 38060 82016 38124 82080
rect 38140 82016 38204 82080
rect 38220 82016 38284 82080
rect 43740 82016 43804 82080
rect 43820 82016 43884 82080
rect 43900 82016 43964 82080
rect 43980 82016 44044 82080
rect 44060 82016 44124 82080
rect 44140 82016 44204 82080
rect 44220 82016 44284 82080
rect 49740 82076 49804 82080
rect 49740 82020 49742 82076
rect 49742 82020 49798 82076
rect 49798 82020 49804 82076
rect 49740 82016 49804 82020
rect 49820 82016 49884 82080
rect 49900 82016 49964 82080
rect 49980 82016 50044 82080
rect 50060 82016 50124 82080
rect 50140 82016 50204 82080
rect 50220 82016 50284 82080
rect 55740 82016 55804 82080
rect 55820 82016 55884 82080
rect 55900 82016 55964 82080
rect 55980 82016 56044 82080
rect 56060 82016 56124 82080
rect 56140 82016 56204 82080
rect 56220 82016 56284 82080
rect 61740 82016 61804 82080
rect 61820 82016 61884 82080
rect 61900 82016 61964 82080
rect 61980 82016 62044 82080
rect 62060 82016 62124 82080
rect 62140 82016 62204 82080
rect 62220 82016 62284 82080
rect 67740 82016 67804 82080
rect 67820 82016 67884 82080
rect 67900 82016 67964 82080
rect 67980 82016 68044 82080
rect 68060 82016 68124 82080
rect 68140 82016 68204 82080
rect 68220 82016 68284 82080
rect 73740 82016 73804 82080
rect 73820 82016 73884 82080
rect 73900 82016 73964 82080
rect 73980 82016 74044 82080
rect 74060 82016 74124 82080
rect 74140 82016 74204 82080
rect 74220 82016 74284 82080
rect 1740 81936 1804 82000
rect 1820 81936 1884 82000
rect 1900 81936 1964 82000
rect 1980 81936 2044 82000
rect 2060 81936 2124 82000
rect 2140 81996 2204 82000
rect 2220 81996 2284 82000
rect 2140 81940 2184 81996
rect 2184 81940 2204 81996
rect 2220 81940 2240 81996
rect 2240 81940 2264 81996
rect 2264 81940 2284 81996
rect 2140 81936 2204 81940
rect 2220 81936 2284 81940
rect 7740 81936 7804 82000
rect 7820 81936 7884 82000
rect 7900 81936 7964 82000
rect 7980 81936 8044 82000
rect 8060 81936 8124 82000
rect 8140 81936 8204 82000
rect 8220 81996 8284 82000
rect 8220 81940 8283 81996
rect 8283 81940 8284 81996
rect 8220 81936 8284 81940
rect 13740 81936 13804 82000
rect 13820 81936 13884 82000
rect 13900 81936 13964 82000
rect 13980 81936 14044 82000
rect 14060 81996 14124 82000
rect 14060 81940 14063 81996
rect 14063 81940 14119 81996
rect 14119 81940 14124 81996
rect 14060 81936 14124 81940
rect 14140 81936 14204 82000
rect 14220 81936 14284 82000
rect 19740 81936 19804 82000
rect 19820 81996 19884 82000
rect 19820 81940 19843 81996
rect 19843 81940 19884 81996
rect 19820 81936 19884 81940
rect 19900 81936 19964 82000
rect 19980 81936 20044 82000
rect 20060 81936 20124 82000
rect 20140 81936 20204 82000
rect 20220 81936 20284 82000
rect 25740 81936 25804 82000
rect 25820 81936 25884 82000
rect 25900 81936 25964 82000
rect 25980 81936 26044 82000
rect 26060 81936 26124 82000
rect 26140 81936 26204 82000
rect 26220 81936 26284 82000
rect 31740 81936 31804 82000
rect 31820 81936 31884 82000
rect 31900 81936 31964 82000
rect 31980 81936 32044 82000
rect 32060 81936 32124 82000
rect 32140 81936 32204 82000
rect 32220 81936 32284 82000
rect 37740 81936 37804 82000
rect 37820 81936 37884 82000
rect 37900 81936 37964 82000
rect 37980 81936 38044 82000
rect 38060 81936 38124 82000
rect 38140 81936 38204 82000
rect 38220 81936 38284 82000
rect 43740 81936 43804 82000
rect 43820 81936 43884 82000
rect 43900 81936 43964 82000
rect 43980 81936 44044 82000
rect 44060 81936 44124 82000
rect 44140 81936 44204 82000
rect 44220 81936 44284 82000
rect 49740 81996 49804 82000
rect 49740 81940 49742 81996
rect 49742 81940 49798 81996
rect 49798 81940 49804 81996
rect 49740 81936 49804 81940
rect 49820 81936 49884 82000
rect 49900 81936 49964 82000
rect 49980 81936 50044 82000
rect 50060 81936 50124 82000
rect 50140 81936 50204 82000
rect 50220 81936 50284 82000
rect 55740 81936 55804 82000
rect 55820 81936 55884 82000
rect 55900 81936 55964 82000
rect 55980 81936 56044 82000
rect 56060 81936 56124 82000
rect 56140 81936 56204 82000
rect 56220 81936 56284 82000
rect 61740 81936 61804 82000
rect 61820 81936 61884 82000
rect 61900 81936 61964 82000
rect 61980 81936 62044 82000
rect 62060 81936 62124 82000
rect 62140 81936 62204 82000
rect 62220 81936 62284 82000
rect 67740 81936 67804 82000
rect 67820 81936 67884 82000
rect 67900 81936 67964 82000
rect 67980 81936 68044 82000
rect 68060 81936 68124 82000
rect 68140 81936 68204 82000
rect 68220 81936 68284 82000
rect 73740 81936 73804 82000
rect 73820 81936 73884 82000
rect 73900 81936 73964 82000
rect 73980 81936 74044 82000
rect 74060 81936 74124 82000
rect 74140 81936 74204 82000
rect 74220 81936 74284 82000
rect 4740 74528 4804 74592
rect 4820 74528 4884 74592
rect 4900 74528 4964 74592
rect 4980 74528 5044 74592
rect 5060 74528 5124 74592
rect 5140 74528 5204 74592
rect 5220 74528 5284 74592
rect 10740 74528 10804 74592
rect 10820 74528 10884 74592
rect 10900 74528 10964 74592
rect 10980 74528 11044 74592
rect 11060 74528 11124 74592
rect 11140 74528 11204 74592
rect 11220 74528 11284 74592
rect 16740 74528 16804 74592
rect 16820 74528 16884 74592
rect 16900 74528 16964 74592
rect 16980 74528 17044 74592
rect 17060 74588 17124 74592
rect 17140 74588 17204 74592
rect 17060 74532 17100 74588
rect 17100 74532 17124 74588
rect 17140 74532 17156 74588
rect 17156 74532 17204 74588
rect 17060 74528 17124 74532
rect 17140 74528 17204 74532
rect 17220 74528 17284 74592
rect 22740 74528 22804 74592
rect 22820 74588 22884 74592
rect 22900 74588 22964 74592
rect 22820 74532 22880 74588
rect 22880 74532 22884 74588
rect 22900 74532 22936 74588
rect 22936 74532 22964 74588
rect 22820 74528 22884 74532
rect 22900 74528 22964 74532
rect 22980 74528 23044 74592
rect 23060 74528 23124 74592
rect 23140 74528 23204 74592
rect 23220 74528 23284 74592
rect 28740 74528 28804 74592
rect 28820 74528 28884 74592
rect 28900 74528 28964 74592
rect 28980 74528 29044 74592
rect 29060 74528 29124 74592
rect 29140 74528 29204 74592
rect 29220 74528 29284 74592
rect 34740 74528 34804 74592
rect 34820 74528 34884 74592
rect 34900 74528 34964 74592
rect 34980 74528 35044 74592
rect 35060 74528 35124 74592
rect 35140 74528 35204 74592
rect 35220 74528 35284 74592
rect 40740 74528 40804 74592
rect 40820 74528 40884 74592
rect 40900 74528 40964 74592
rect 40980 74528 41044 74592
rect 41060 74528 41124 74592
rect 41140 74528 41204 74592
rect 41220 74528 41284 74592
rect 46740 74528 46804 74592
rect 46820 74528 46884 74592
rect 46900 74528 46964 74592
rect 46980 74528 47044 74592
rect 47060 74528 47124 74592
rect 47140 74528 47204 74592
rect 47220 74528 47284 74592
rect 52740 74528 52804 74592
rect 52820 74528 52884 74592
rect 52900 74528 52964 74592
rect 52980 74528 53044 74592
rect 53060 74528 53124 74592
rect 53140 74528 53204 74592
rect 53220 74528 53284 74592
rect 58740 74528 58804 74592
rect 58820 74528 58884 74592
rect 58900 74528 58964 74592
rect 58980 74528 59044 74592
rect 59060 74588 59124 74592
rect 59060 74532 59104 74588
rect 59104 74532 59124 74588
rect 59060 74528 59124 74532
rect 59140 74528 59204 74592
rect 59220 74528 59284 74592
rect 64740 74528 64804 74592
rect 64820 74528 64884 74592
rect 64900 74528 64964 74592
rect 64980 74528 65044 74592
rect 65060 74528 65124 74592
rect 65140 74528 65204 74592
rect 65220 74528 65284 74592
rect 70740 74528 70804 74592
rect 70820 74528 70884 74592
rect 70900 74528 70964 74592
rect 70980 74528 71044 74592
rect 71060 74528 71124 74592
rect 71140 74528 71204 74592
rect 71220 74528 71284 74592
rect 4740 74448 4804 74512
rect 4820 74448 4884 74512
rect 4900 74448 4964 74512
rect 4980 74448 5044 74512
rect 5060 74448 5124 74512
rect 5140 74448 5204 74512
rect 5220 74448 5284 74512
rect 10740 74448 10804 74512
rect 10820 74448 10884 74512
rect 10900 74448 10964 74512
rect 10980 74448 11044 74512
rect 11060 74448 11124 74512
rect 11140 74448 11204 74512
rect 11220 74448 11284 74512
rect 16740 74448 16804 74512
rect 16820 74448 16884 74512
rect 16900 74448 16964 74512
rect 16980 74448 17044 74512
rect 17060 74508 17124 74512
rect 17140 74508 17204 74512
rect 17060 74452 17100 74508
rect 17100 74452 17124 74508
rect 17140 74452 17156 74508
rect 17156 74452 17204 74508
rect 17060 74448 17124 74452
rect 17140 74448 17204 74452
rect 17220 74448 17284 74512
rect 22740 74448 22804 74512
rect 22820 74508 22884 74512
rect 22900 74508 22964 74512
rect 22820 74452 22880 74508
rect 22880 74452 22884 74508
rect 22900 74452 22936 74508
rect 22936 74452 22964 74508
rect 22820 74448 22884 74452
rect 22900 74448 22964 74452
rect 22980 74448 23044 74512
rect 23060 74448 23124 74512
rect 23140 74448 23204 74512
rect 23220 74448 23284 74512
rect 28740 74448 28804 74512
rect 28820 74448 28884 74512
rect 28900 74448 28964 74512
rect 28980 74448 29044 74512
rect 29060 74448 29124 74512
rect 29140 74448 29204 74512
rect 29220 74448 29284 74512
rect 34740 74448 34804 74512
rect 34820 74448 34884 74512
rect 34900 74448 34964 74512
rect 34980 74448 35044 74512
rect 35060 74448 35124 74512
rect 35140 74448 35204 74512
rect 35220 74448 35284 74512
rect 40740 74448 40804 74512
rect 40820 74448 40884 74512
rect 40900 74448 40964 74512
rect 40980 74448 41044 74512
rect 41060 74448 41124 74512
rect 41140 74448 41204 74512
rect 41220 74448 41284 74512
rect 46740 74448 46804 74512
rect 46820 74448 46884 74512
rect 46900 74448 46964 74512
rect 46980 74448 47044 74512
rect 47060 74448 47124 74512
rect 47140 74448 47204 74512
rect 47220 74448 47284 74512
rect 52740 74448 52804 74512
rect 52820 74448 52884 74512
rect 52900 74448 52964 74512
rect 52980 74448 53044 74512
rect 53060 74448 53124 74512
rect 53140 74448 53204 74512
rect 53220 74448 53284 74512
rect 58740 74448 58804 74512
rect 58820 74448 58884 74512
rect 58900 74448 58964 74512
rect 58980 74448 59044 74512
rect 59060 74508 59124 74512
rect 59060 74452 59104 74508
rect 59104 74452 59124 74508
rect 59060 74448 59124 74452
rect 59140 74448 59204 74512
rect 59220 74448 59284 74512
rect 64740 74448 64804 74512
rect 64820 74448 64884 74512
rect 64900 74448 64964 74512
rect 64980 74448 65044 74512
rect 65060 74448 65124 74512
rect 65140 74448 65204 74512
rect 65220 74448 65284 74512
rect 70740 74448 70804 74512
rect 70820 74448 70884 74512
rect 70900 74448 70964 74512
rect 70980 74448 71044 74512
rect 71060 74448 71124 74512
rect 71140 74448 71204 74512
rect 71220 74448 71284 74512
rect 4740 74368 4804 74432
rect 4820 74368 4884 74432
rect 4900 74368 4964 74432
rect 4980 74368 5044 74432
rect 5060 74368 5124 74432
rect 5140 74368 5204 74432
rect 5220 74368 5284 74432
rect 10740 74368 10804 74432
rect 10820 74368 10884 74432
rect 10900 74368 10964 74432
rect 10980 74368 11044 74432
rect 11060 74368 11124 74432
rect 11140 74368 11204 74432
rect 11220 74368 11284 74432
rect 16740 74368 16804 74432
rect 16820 74368 16884 74432
rect 16900 74368 16964 74432
rect 16980 74368 17044 74432
rect 17060 74428 17124 74432
rect 17140 74428 17204 74432
rect 17060 74372 17100 74428
rect 17100 74372 17124 74428
rect 17140 74372 17156 74428
rect 17156 74372 17204 74428
rect 17060 74368 17124 74372
rect 17140 74368 17204 74372
rect 17220 74368 17284 74432
rect 22740 74368 22804 74432
rect 22820 74428 22884 74432
rect 22900 74428 22964 74432
rect 22820 74372 22880 74428
rect 22880 74372 22884 74428
rect 22900 74372 22936 74428
rect 22936 74372 22964 74428
rect 22820 74368 22884 74372
rect 22900 74368 22964 74372
rect 22980 74368 23044 74432
rect 23060 74368 23124 74432
rect 23140 74368 23204 74432
rect 23220 74368 23284 74432
rect 28740 74368 28804 74432
rect 28820 74368 28884 74432
rect 28900 74368 28964 74432
rect 28980 74368 29044 74432
rect 29060 74368 29124 74432
rect 29140 74368 29204 74432
rect 29220 74368 29284 74432
rect 34740 74368 34804 74432
rect 34820 74368 34884 74432
rect 34900 74368 34964 74432
rect 34980 74368 35044 74432
rect 35060 74368 35124 74432
rect 35140 74368 35204 74432
rect 35220 74368 35284 74432
rect 40740 74368 40804 74432
rect 40820 74368 40884 74432
rect 40900 74368 40964 74432
rect 40980 74368 41044 74432
rect 41060 74368 41124 74432
rect 41140 74368 41204 74432
rect 41220 74368 41284 74432
rect 46740 74368 46804 74432
rect 46820 74368 46884 74432
rect 46900 74368 46964 74432
rect 46980 74368 47044 74432
rect 47060 74368 47124 74432
rect 47140 74368 47204 74432
rect 47220 74368 47284 74432
rect 52740 74368 52804 74432
rect 52820 74368 52884 74432
rect 52900 74368 52964 74432
rect 52980 74368 53044 74432
rect 53060 74368 53124 74432
rect 53140 74368 53204 74432
rect 53220 74368 53284 74432
rect 58740 74368 58804 74432
rect 58820 74368 58884 74432
rect 58900 74368 58964 74432
rect 58980 74368 59044 74432
rect 59060 74428 59124 74432
rect 59060 74372 59104 74428
rect 59104 74372 59124 74428
rect 59060 74368 59124 74372
rect 59140 74368 59204 74432
rect 59220 74368 59284 74432
rect 64740 74368 64804 74432
rect 64820 74368 64884 74432
rect 64900 74368 64964 74432
rect 64980 74368 65044 74432
rect 65060 74368 65124 74432
rect 65140 74368 65204 74432
rect 65220 74368 65284 74432
rect 70740 74368 70804 74432
rect 70820 74368 70884 74432
rect 70900 74368 70964 74432
rect 70980 74368 71044 74432
rect 71060 74368 71124 74432
rect 71140 74368 71204 74432
rect 71220 74368 71284 74432
rect 4740 74288 4804 74352
rect 4820 74288 4884 74352
rect 4900 74288 4964 74352
rect 4980 74288 5044 74352
rect 5060 74288 5124 74352
rect 5140 74288 5204 74352
rect 5220 74288 5284 74352
rect 10740 74288 10804 74352
rect 10820 74288 10884 74352
rect 10900 74288 10964 74352
rect 10980 74288 11044 74352
rect 11060 74288 11124 74352
rect 11140 74288 11204 74352
rect 11220 74288 11284 74352
rect 16740 74288 16804 74352
rect 16820 74288 16884 74352
rect 16900 74288 16964 74352
rect 16980 74288 17044 74352
rect 17060 74348 17124 74352
rect 17140 74348 17204 74352
rect 17060 74292 17100 74348
rect 17100 74292 17124 74348
rect 17140 74292 17156 74348
rect 17156 74292 17204 74348
rect 17060 74288 17124 74292
rect 17140 74288 17204 74292
rect 17220 74288 17284 74352
rect 22740 74288 22804 74352
rect 22820 74348 22884 74352
rect 22900 74348 22964 74352
rect 22820 74292 22880 74348
rect 22880 74292 22884 74348
rect 22900 74292 22936 74348
rect 22936 74292 22964 74348
rect 22820 74288 22884 74292
rect 22900 74288 22964 74292
rect 22980 74288 23044 74352
rect 23060 74288 23124 74352
rect 23140 74288 23204 74352
rect 23220 74288 23284 74352
rect 28740 74288 28804 74352
rect 28820 74288 28884 74352
rect 28900 74288 28964 74352
rect 28980 74288 29044 74352
rect 29060 74288 29124 74352
rect 29140 74288 29204 74352
rect 29220 74288 29284 74352
rect 34740 74288 34804 74352
rect 34820 74288 34884 74352
rect 34900 74288 34964 74352
rect 34980 74288 35044 74352
rect 35060 74288 35124 74352
rect 35140 74288 35204 74352
rect 35220 74288 35284 74352
rect 40740 74288 40804 74352
rect 40820 74288 40884 74352
rect 40900 74288 40964 74352
rect 40980 74288 41044 74352
rect 41060 74288 41124 74352
rect 41140 74288 41204 74352
rect 41220 74288 41284 74352
rect 46740 74288 46804 74352
rect 46820 74288 46884 74352
rect 46900 74288 46964 74352
rect 46980 74288 47044 74352
rect 47060 74288 47124 74352
rect 47140 74288 47204 74352
rect 47220 74288 47284 74352
rect 52740 74288 52804 74352
rect 52820 74288 52884 74352
rect 52900 74288 52964 74352
rect 52980 74288 53044 74352
rect 53060 74288 53124 74352
rect 53140 74288 53204 74352
rect 53220 74288 53284 74352
rect 58740 74288 58804 74352
rect 58820 74288 58884 74352
rect 58900 74288 58964 74352
rect 58980 74288 59044 74352
rect 59060 74348 59124 74352
rect 59060 74292 59104 74348
rect 59104 74292 59124 74348
rect 59060 74288 59124 74292
rect 59140 74288 59204 74352
rect 59220 74288 59284 74352
rect 64740 74288 64804 74352
rect 64820 74288 64884 74352
rect 64900 74288 64964 74352
rect 64980 74288 65044 74352
rect 65060 74288 65124 74352
rect 65140 74288 65204 74352
rect 65220 74288 65284 74352
rect 70740 74288 70804 74352
rect 70820 74288 70884 74352
rect 70900 74288 70964 74352
rect 70980 74288 71044 74352
rect 71060 74288 71124 74352
rect 71140 74288 71204 74352
rect 71220 74288 71284 74352
rect 1740 72176 1804 72240
rect 1820 72176 1884 72240
rect 1900 72176 1964 72240
rect 1980 72176 2044 72240
rect 2060 72176 2124 72240
rect 2140 72236 2204 72240
rect 2220 72236 2284 72240
rect 2140 72180 2184 72236
rect 2184 72180 2204 72236
rect 2220 72180 2240 72236
rect 2240 72180 2264 72236
rect 2264 72180 2284 72236
rect 2140 72176 2204 72180
rect 2220 72176 2284 72180
rect 7740 72176 7804 72240
rect 7820 72176 7884 72240
rect 7900 72176 7964 72240
rect 7980 72176 8044 72240
rect 8060 72176 8124 72240
rect 8140 72176 8204 72240
rect 8220 72236 8284 72240
rect 8220 72180 8283 72236
rect 8283 72180 8284 72236
rect 8220 72176 8284 72180
rect 13740 72176 13804 72240
rect 13820 72176 13884 72240
rect 13900 72176 13964 72240
rect 13980 72176 14044 72240
rect 14060 72236 14124 72240
rect 14060 72180 14063 72236
rect 14063 72180 14119 72236
rect 14119 72180 14124 72236
rect 14060 72176 14124 72180
rect 14140 72176 14204 72240
rect 14220 72176 14284 72240
rect 19740 72176 19804 72240
rect 19820 72236 19884 72240
rect 19820 72180 19843 72236
rect 19843 72180 19884 72236
rect 19820 72176 19884 72180
rect 19900 72176 19964 72240
rect 19980 72176 20044 72240
rect 20060 72176 20124 72240
rect 20140 72176 20204 72240
rect 20220 72176 20284 72240
rect 25740 72176 25804 72240
rect 25820 72176 25884 72240
rect 25900 72176 25964 72240
rect 25980 72176 26044 72240
rect 26060 72176 26124 72240
rect 26140 72176 26204 72240
rect 26220 72176 26284 72240
rect 31740 72176 31804 72240
rect 31820 72176 31884 72240
rect 31900 72176 31964 72240
rect 31980 72176 32044 72240
rect 32060 72176 32124 72240
rect 32140 72176 32204 72240
rect 32220 72176 32284 72240
rect 37740 72176 37804 72240
rect 37820 72176 37884 72240
rect 37900 72176 37964 72240
rect 37980 72176 38044 72240
rect 38060 72176 38124 72240
rect 38140 72176 38204 72240
rect 38220 72176 38284 72240
rect 43740 72176 43804 72240
rect 43820 72176 43884 72240
rect 43900 72176 43964 72240
rect 43980 72176 44044 72240
rect 44060 72176 44124 72240
rect 44140 72176 44204 72240
rect 44220 72176 44284 72240
rect 49740 72236 49804 72240
rect 49740 72180 49742 72236
rect 49742 72180 49798 72236
rect 49798 72180 49804 72236
rect 49740 72176 49804 72180
rect 49820 72176 49884 72240
rect 49900 72176 49964 72240
rect 49980 72176 50044 72240
rect 50060 72176 50124 72240
rect 50140 72176 50204 72240
rect 50220 72176 50284 72240
rect 55740 72176 55804 72240
rect 55820 72176 55884 72240
rect 55900 72176 55964 72240
rect 55980 72176 56044 72240
rect 56060 72176 56124 72240
rect 56140 72176 56204 72240
rect 56220 72176 56284 72240
rect 61740 72176 61804 72240
rect 61820 72176 61884 72240
rect 61900 72176 61964 72240
rect 61980 72176 62044 72240
rect 62060 72176 62124 72240
rect 62140 72176 62204 72240
rect 62220 72176 62284 72240
rect 67740 72176 67804 72240
rect 67820 72176 67884 72240
rect 67900 72176 67964 72240
rect 67980 72176 68044 72240
rect 68060 72176 68124 72240
rect 68140 72176 68204 72240
rect 68220 72176 68284 72240
rect 73740 72176 73804 72240
rect 73820 72176 73884 72240
rect 73900 72176 73964 72240
rect 73980 72176 74044 72240
rect 74060 72176 74124 72240
rect 74140 72176 74204 72240
rect 74220 72176 74284 72240
rect 1740 72096 1804 72160
rect 1820 72096 1884 72160
rect 1900 72096 1964 72160
rect 1980 72096 2044 72160
rect 2060 72096 2124 72160
rect 2140 72156 2204 72160
rect 2220 72156 2284 72160
rect 2140 72100 2184 72156
rect 2184 72100 2204 72156
rect 2220 72100 2240 72156
rect 2240 72100 2264 72156
rect 2264 72100 2284 72156
rect 2140 72096 2204 72100
rect 2220 72096 2284 72100
rect 7740 72096 7804 72160
rect 7820 72096 7884 72160
rect 7900 72096 7964 72160
rect 7980 72096 8044 72160
rect 8060 72096 8124 72160
rect 8140 72096 8204 72160
rect 8220 72156 8284 72160
rect 8220 72100 8283 72156
rect 8283 72100 8284 72156
rect 8220 72096 8284 72100
rect 13740 72096 13804 72160
rect 13820 72096 13884 72160
rect 13900 72096 13964 72160
rect 13980 72096 14044 72160
rect 14060 72156 14124 72160
rect 14060 72100 14063 72156
rect 14063 72100 14119 72156
rect 14119 72100 14124 72156
rect 14060 72096 14124 72100
rect 14140 72096 14204 72160
rect 14220 72096 14284 72160
rect 19740 72096 19804 72160
rect 19820 72156 19884 72160
rect 19820 72100 19843 72156
rect 19843 72100 19884 72156
rect 19820 72096 19884 72100
rect 19900 72096 19964 72160
rect 19980 72096 20044 72160
rect 20060 72096 20124 72160
rect 20140 72096 20204 72160
rect 20220 72096 20284 72160
rect 25740 72096 25804 72160
rect 25820 72096 25884 72160
rect 25900 72096 25964 72160
rect 25980 72096 26044 72160
rect 26060 72096 26124 72160
rect 26140 72096 26204 72160
rect 26220 72096 26284 72160
rect 31740 72096 31804 72160
rect 31820 72096 31884 72160
rect 31900 72096 31964 72160
rect 31980 72096 32044 72160
rect 32060 72096 32124 72160
rect 32140 72096 32204 72160
rect 32220 72096 32284 72160
rect 37740 72096 37804 72160
rect 37820 72096 37884 72160
rect 37900 72096 37964 72160
rect 37980 72096 38044 72160
rect 38060 72096 38124 72160
rect 38140 72096 38204 72160
rect 38220 72096 38284 72160
rect 43740 72096 43804 72160
rect 43820 72096 43884 72160
rect 43900 72096 43964 72160
rect 43980 72096 44044 72160
rect 44060 72096 44124 72160
rect 44140 72096 44204 72160
rect 44220 72096 44284 72160
rect 49740 72156 49804 72160
rect 49740 72100 49742 72156
rect 49742 72100 49798 72156
rect 49798 72100 49804 72156
rect 49740 72096 49804 72100
rect 49820 72096 49884 72160
rect 49900 72096 49964 72160
rect 49980 72096 50044 72160
rect 50060 72096 50124 72160
rect 50140 72096 50204 72160
rect 50220 72096 50284 72160
rect 55740 72096 55804 72160
rect 55820 72096 55884 72160
rect 55900 72096 55964 72160
rect 55980 72096 56044 72160
rect 56060 72096 56124 72160
rect 56140 72096 56204 72160
rect 56220 72096 56284 72160
rect 61740 72096 61804 72160
rect 61820 72096 61884 72160
rect 61900 72096 61964 72160
rect 61980 72096 62044 72160
rect 62060 72096 62124 72160
rect 62140 72096 62204 72160
rect 62220 72096 62284 72160
rect 67740 72096 67804 72160
rect 67820 72096 67884 72160
rect 67900 72096 67964 72160
rect 67980 72096 68044 72160
rect 68060 72096 68124 72160
rect 68140 72096 68204 72160
rect 68220 72096 68284 72160
rect 73740 72096 73804 72160
rect 73820 72096 73884 72160
rect 73900 72096 73964 72160
rect 73980 72096 74044 72160
rect 74060 72096 74124 72160
rect 74140 72096 74204 72160
rect 74220 72096 74284 72160
rect 1740 72016 1804 72080
rect 1820 72016 1884 72080
rect 1900 72016 1964 72080
rect 1980 72016 2044 72080
rect 2060 72016 2124 72080
rect 2140 72076 2204 72080
rect 2220 72076 2284 72080
rect 2140 72020 2184 72076
rect 2184 72020 2204 72076
rect 2220 72020 2240 72076
rect 2240 72020 2264 72076
rect 2264 72020 2284 72076
rect 2140 72016 2204 72020
rect 2220 72016 2284 72020
rect 7740 72016 7804 72080
rect 7820 72016 7884 72080
rect 7900 72016 7964 72080
rect 7980 72016 8044 72080
rect 8060 72016 8124 72080
rect 8140 72016 8204 72080
rect 8220 72076 8284 72080
rect 8220 72020 8283 72076
rect 8283 72020 8284 72076
rect 8220 72016 8284 72020
rect 13740 72016 13804 72080
rect 13820 72016 13884 72080
rect 13900 72016 13964 72080
rect 13980 72016 14044 72080
rect 14060 72076 14124 72080
rect 14060 72020 14063 72076
rect 14063 72020 14119 72076
rect 14119 72020 14124 72076
rect 14060 72016 14124 72020
rect 14140 72016 14204 72080
rect 14220 72016 14284 72080
rect 19740 72016 19804 72080
rect 19820 72076 19884 72080
rect 19820 72020 19843 72076
rect 19843 72020 19884 72076
rect 19820 72016 19884 72020
rect 19900 72016 19964 72080
rect 19980 72016 20044 72080
rect 20060 72016 20124 72080
rect 20140 72016 20204 72080
rect 20220 72016 20284 72080
rect 25740 72016 25804 72080
rect 25820 72016 25884 72080
rect 25900 72016 25964 72080
rect 25980 72016 26044 72080
rect 26060 72016 26124 72080
rect 26140 72016 26204 72080
rect 26220 72016 26284 72080
rect 31740 72016 31804 72080
rect 31820 72016 31884 72080
rect 31900 72016 31964 72080
rect 31980 72016 32044 72080
rect 32060 72016 32124 72080
rect 32140 72016 32204 72080
rect 32220 72016 32284 72080
rect 37740 72016 37804 72080
rect 37820 72016 37884 72080
rect 37900 72016 37964 72080
rect 37980 72016 38044 72080
rect 38060 72016 38124 72080
rect 38140 72016 38204 72080
rect 38220 72016 38284 72080
rect 43740 72016 43804 72080
rect 43820 72016 43884 72080
rect 43900 72016 43964 72080
rect 43980 72016 44044 72080
rect 44060 72016 44124 72080
rect 44140 72016 44204 72080
rect 44220 72016 44284 72080
rect 49740 72076 49804 72080
rect 49740 72020 49742 72076
rect 49742 72020 49798 72076
rect 49798 72020 49804 72076
rect 49740 72016 49804 72020
rect 49820 72016 49884 72080
rect 49900 72016 49964 72080
rect 49980 72016 50044 72080
rect 50060 72016 50124 72080
rect 50140 72016 50204 72080
rect 50220 72016 50284 72080
rect 55740 72016 55804 72080
rect 55820 72016 55884 72080
rect 55900 72016 55964 72080
rect 55980 72016 56044 72080
rect 56060 72016 56124 72080
rect 56140 72016 56204 72080
rect 56220 72016 56284 72080
rect 61740 72016 61804 72080
rect 61820 72016 61884 72080
rect 61900 72016 61964 72080
rect 61980 72016 62044 72080
rect 62060 72016 62124 72080
rect 62140 72016 62204 72080
rect 62220 72016 62284 72080
rect 67740 72016 67804 72080
rect 67820 72016 67884 72080
rect 67900 72016 67964 72080
rect 67980 72016 68044 72080
rect 68060 72016 68124 72080
rect 68140 72016 68204 72080
rect 68220 72016 68284 72080
rect 73740 72016 73804 72080
rect 73820 72016 73884 72080
rect 73900 72016 73964 72080
rect 73980 72016 74044 72080
rect 74060 72016 74124 72080
rect 74140 72016 74204 72080
rect 74220 72016 74284 72080
rect 1740 71936 1804 72000
rect 1820 71936 1884 72000
rect 1900 71936 1964 72000
rect 1980 71936 2044 72000
rect 2060 71936 2124 72000
rect 2140 71996 2204 72000
rect 2220 71996 2284 72000
rect 2140 71940 2184 71996
rect 2184 71940 2204 71996
rect 2220 71940 2240 71996
rect 2240 71940 2264 71996
rect 2264 71940 2284 71996
rect 2140 71936 2204 71940
rect 2220 71936 2284 71940
rect 7740 71936 7804 72000
rect 7820 71936 7884 72000
rect 7900 71936 7964 72000
rect 7980 71936 8044 72000
rect 8060 71936 8124 72000
rect 8140 71936 8204 72000
rect 8220 71996 8284 72000
rect 8220 71940 8283 71996
rect 8283 71940 8284 71996
rect 8220 71936 8284 71940
rect 13740 71936 13804 72000
rect 13820 71936 13884 72000
rect 13900 71936 13964 72000
rect 13980 71936 14044 72000
rect 14060 71996 14124 72000
rect 14060 71940 14063 71996
rect 14063 71940 14119 71996
rect 14119 71940 14124 71996
rect 14060 71936 14124 71940
rect 14140 71936 14204 72000
rect 14220 71936 14284 72000
rect 19740 71936 19804 72000
rect 19820 71996 19884 72000
rect 19820 71940 19843 71996
rect 19843 71940 19884 71996
rect 19820 71936 19884 71940
rect 19900 71936 19964 72000
rect 19980 71936 20044 72000
rect 20060 71936 20124 72000
rect 20140 71936 20204 72000
rect 20220 71936 20284 72000
rect 25740 71936 25804 72000
rect 25820 71936 25884 72000
rect 25900 71936 25964 72000
rect 25980 71936 26044 72000
rect 26060 71936 26124 72000
rect 26140 71936 26204 72000
rect 26220 71936 26284 72000
rect 31740 71936 31804 72000
rect 31820 71936 31884 72000
rect 31900 71936 31964 72000
rect 31980 71936 32044 72000
rect 32060 71936 32124 72000
rect 32140 71936 32204 72000
rect 32220 71936 32284 72000
rect 37740 71936 37804 72000
rect 37820 71936 37884 72000
rect 37900 71936 37964 72000
rect 37980 71936 38044 72000
rect 38060 71936 38124 72000
rect 38140 71936 38204 72000
rect 38220 71936 38284 72000
rect 43740 71936 43804 72000
rect 43820 71936 43884 72000
rect 43900 71936 43964 72000
rect 43980 71936 44044 72000
rect 44060 71936 44124 72000
rect 44140 71936 44204 72000
rect 44220 71936 44284 72000
rect 49740 71996 49804 72000
rect 49740 71940 49742 71996
rect 49742 71940 49798 71996
rect 49798 71940 49804 71996
rect 49740 71936 49804 71940
rect 49820 71936 49884 72000
rect 49900 71936 49964 72000
rect 49980 71936 50044 72000
rect 50060 71936 50124 72000
rect 50140 71936 50204 72000
rect 50220 71936 50284 72000
rect 55740 71936 55804 72000
rect 55820 71936 55884 72000
rect 55900 71936 55964 72000
rect 55980 71936 56044 72000
rect 56060 71936 56124 72000
rect 56140 71936 56204 72000
rect 56220 71936 56284 72000
rect 61740 71936 61804 72000
rect 61820 71936 61884 72000
rect 61900 71936 61964 72000
rect 61980 71936 62044 72000
rect 62060 71936 62124 72000
rect 62140 71936 62204 72000
rect 62220 71936 62284 72000
rect 67740 71936 67804 72000
rect 67820 71936 67884 72000
rect 67900 71936 67964 72000
rect 67980 71936 68044 72000
rect 68060 71936 68124 72000
rect 68140 71936 68204 72000
rect 68220 71936 68284 72000
rect 73740 71936 73804 72000
rect 73820 71936 73884 72000
rect 73900 71936 73964 72000
rect 73980 71936 74044 72000
rect 74060 71936 74124 72000
rect 74140 71936 74204 72000
rect 74220 71936 74284 72000
rect 4740 64528 4804 64592
rect 4820 64528 4884 64592
rect 4900 64528 4964 64592
rect 4980 64528 5044 64592
rect 5060 64528 5124 64592
rect 5140 64528 5204 64592
rect 5220 64528 5284 64592
rect 10740 64528 10804 64592
rect 10820 64528 10884 64592
rect 10900 64528 10964 64592
rect 10980 64528 11044 64592
rect 11060 64528 11124 64592
rect 11140 64528 11204 64592
rect 11220 64528 11284 64592
rect 16740 64528 16804 64592
rect 16820 64528 16884 64592
rect 16900 64528 16964 64592
rect 16980 64528 17044 64592
rect 17060 64588 17124 64592
rect 17140 64588 17204 64592
rect 17060 64532 17100 64588
rect 17100 64532 17124 64588
rect 17140 64532 17156 64588
rect 17156 64532 17204 64588
rect 17060 64528 17124 64532
rect 17140 64528 17204 64532
rect 17220 64528 17284 64592
rect 22740 64528 22804 64592
rect 22820 64588 22884 64592
rect 22900 64588 22964 64592
rect 22820 64532 22880 64588
rect 22880 64532 22884 64588
rect 22900 64532 22936 64588
rect 22936 64532 22964 64588
rect 22820 64528 22884 64532
rect 22900 64528 22964 64532
rect 22980 64528 23044 64592
rect 23060 64528 23124 64592
rect 23140 64528 23204 64592
rect 23220 64528 23284 64592
rect 28740 64528 28804 64592
rect 28820 64528 28884 64592
rect 28900 64528 28964 64592
rect 28980 64528 29044 64592
rect 29060 64528 29124 64592
rect 29140 64528 29204 64592
rect 29220 64528 29284 64592
rect 34740 64528 34804 64592
rect 34820 64528 34884 64592
rect 34900 64528 34964 64592
rect 34980 64528 35044 64592
rect 35060 64528 35124 64592
rect 35140 64528 35204 64592
rect 35220 64528 35284 64592
rect 40740 64528 40804 64592
rect 40820 64528 40884 64592
rect 40900 64528 40964 64592
rect 40980 64528 41044 64592
rect 41060 64528 41124 64592
rect 41140 64528 41204 64592
rect 41220 64528 41284 64592
rect 46740 64528 46804 64592
rect 46820 64528 46884 64592
rect 46900 64528 46964 64592
rect 46980 64528 47044 64592
rect 47060 64528 47124 64592
rect 47140 64528 47204 64592
rect 47220 64528 47284 64592
rect 52740 64528 52804 64592
rect 52820 64528 52884 64592
rect 52900 64528 52964 64592
rect 52980 64528 53044 64592
rect 53060 64528 53124 64592
rect 53140 64528 53204 64592
rect 53220 64528 53284 64592
rect 58740 64528 58804 64592
rect 58820 64528 58884 64592
rect 58900 64528 58964 64592
rect 58980 64528 59044 64592
rect 59060 64588 59124 64592
rect 59060 64532 59104 64588
rect 59104 64532 59124 64588
rect 59060 64528 59124 64532
rect 59140 64528 59204 64592
rect 59220 64528 59284 64592
rect 64740 64528 64804 64592
rect 64820 64528 64884 64592
rect 64900 64528 64964 64592
rect 64980 64528 65044 64592
rect 65060 64528 65124 64592
rect 65140 64528 65204 64592
rect 65220 64528 65284 64592
rect 70740 64528 70804 64592
rect 70820 64528 70884 64592
rect 70900 64528 70964 64592
rect 70980 64528 71044 64592
rect 71060 64528 71124 64592
rect 71140 64528 71204 64592
rect 71220 64528 71284 64592
rect 4740 64448 4804 64512
rect 4820 64448 4884 64512
rect 4900 64448 4964 64512
rect 4980 64448 5044 64512
rect 5060 64448 5124 64512
rect 5140 64448 5204 64512
rect 5220 64448 5284 64512
rect 10740 64448 10804 64512
rect 10820 64448 10884 64512
rect 10900 64448 10964 64512
rect 10980 64448 11044 64512
rect 11060 64448 11124 64512
rect 11140 64448 11204 64512
rect 11220 64448 11284 64512
rect 16740 64448 16804 64512
rect 16820 64448 16884 64512
rect 16900 64448 16964 64512
rect 16980 64448 17044 64512
rect 17060 64508 17124 64512
rect 17140 64508 17204 64512
rect 17060 64452 17100 64508
rect 17100 64452 17124 64508
rect 17140 64452 17156 64508
rect 17156 64452 17204 64508
rect 17060 64448 17124 64452
rect 17140 64448 17204 64452
rect 17220 64448 17284 64512
rect 22740 64448 22804 64512
rect 22820 64508 22884 64512
rect 22900 64508 22964 64512
rect 22820 64452 22880 64508
rect 22880 64452 22884 64508
rect 22900 64452 22936 64508
rect 22936 64452 22964 64508
rect 22820 64448 22884 64452
rect 22900 64448 22964 64452
rect 22980 64448 23044 64512
rect 23060 64448 23124 64512
rect 23140 64448 23204 64512
rect 23220 64448 23284 64512
rect 28740 64448 28804 64512
rect 28820 64448 28884 64512
rect 28900 64448 28964 64512
rect 28980 64448 29044 64512
rect 29060 64448 29124 64512
rect 29140 64448 29204 64512
rect 29220 64448 29284 64512
rect 34740 64448 34804 64512
rect 34820 64448 34884 64512
rect 34900 64448 34964 64512
rect 34980 64448 35044 64512
rect 35060 64448 35124 64512
rect 35140 64448 35204 64512
rect 35220 64448 35284 64512
rect 40740 64448 40804 64512
rect 40820 64448 40884 64512
rect 40900 64448 40964 64512
rect 40980 64448 41044 64512
rect 41060 64448 41124 64512
rect 41140 64448 41204 64512
rect 41220 64448 41284 64512
rect 46740 64448 46804 64512
rect 46820 64448 46884 64512
rect 46900 64448 46964 64512
rect 46980 64448 47044 64512
rect 47060 64448 47124 64512
rect 47140 64448 47204 64512
rect 47220 64448 47284 64512
rect 52740 64448 52804 64512
rect 52820 64448 52884 64512
rect 52900 64448 52964 64512
rect 52980 64448 53044 64512
rect 53060 64448 53124 64512
rect 53140 64448 53204 64512
rect 53220 64448 53284 64512
rect 58740 64448 58804 64512
rect 58820 64448 58884 64512
rect 58900 64448 58964 64512
rect 58980 64448 59044 64512
rect 59060 64508 59124 64512
rect 59060 64452 59104 64508
rect 59104 64452 59124 64508
rect 59060 64448 59124 64452
rect 59140 64448 59204 64512
rect 59220 64448 59284 64512
rect 64740 64448 64804 64512
rect 64820 64448 64884 64512
rect 64900 64448 64964 64512
rect 64980 64448 65044 64512
rect 65060 64448 65124 64512
rect 65140 64448 65204 64512
rect 65220 64448 65284 64512
rect 70740 64448 70804 64512
rect 70820 64448 70884 64512
rect 70900 64448 70964 64512
rect 70980 64448 71044 64512
rect 71060 64448 71124 64512
rect 71140 64448 71204 64512
rect 71220 64448 71284 64512
rect 4740 64368 4804 64432
rect 4820 64368 4884 64432
rect 4900 64368 4964 64432
rect 4980 64368 5044 64432
rect 5060 64368 5124 64432
rect 5140 64368 5204 64432
rect 5220 64368 5284 64432
rect 10740 64368 10804 64432
rect 10820 64368 10884 64432
rect 10900 64368 10964 64432
rect 10980 64368 11044 64432
rect 11060 64368 11124 64432
rect 11140 64368 11204 64432
rect 11220 64368 11284 64432
rect 16740 64368 16804 64432
rect 16820 64368 16884 64432
rect 16900 64368 16964 64432
rect 16980 64368 17044 64432
rect 17060 64428 17124 64432
rect 17140 64428 17204 64432
rect 17060 64372 17100 64428
rect 17100 64372 17124 64428
rect 17140 64372 17156 64428
rect 17156 64372 17204 64428
rect 17060 64368 17124 64372
rect 17140 64368 17204 64372
rect 17220 64368 17284 64432
rect 22740 64368 22804 64432
rect 22820 64428 22884 64432
rect 22900 64428 22964 64432
rect 22820 64372 22880 64428
rect 22880 64372 22884 64428
rect 22900 64372 22936 64428
rect 22936 64372 22964 64428
rect 22820 64368 22884 64372
rect 22900 64368 22964 64372
rect 22980 64368 23044 64432
rect 23060 64368 23124 64432
rect 23140 64368 23204 64432
rect 23220 64368 23284 64432
rect 28740 64368 28804 64432
rect 28820 64368 28884 64432
rect 28900 64368 28964 64432
rect 28980 64368 29044 64432
rect 29060 64368 29124 64432
rect 29140 64368 29204 64432
rect 29220 64368 29284 64432
rect 34740 64368 34804 64432
rect 34820 64368 34884 64432
rect 34900 64368 34964 64432
rect 34980 64368 35044 64432
rect 35060 64368 35124 64432
rect 35140 64368 35204 64432
rect 35220 64368 35284 64432
rect 40740 64368 40804 64432
rect 40820 64368 40884 64432
rect 40900 64368 40964 64432
rect 40980 64368 41044 64432
rect 41060 64368 41124 64432
rect 41140 64368 41204 64432
rect 41220 64368 41284 64432
rect 46740 64368 46804 64432
rect 46820 64368 46884 64432
rect 46900 64368 46964 64432
rect 46980 64368 47044 64432
rect 47060 64368 47124 64432
rect 47140 64368 47204 64432
rect 47220 64368 47284 64432
rect 52740 64368 52804 64432
rect 52820 64368 52884 64432
rect 52900 64368 52964 64432
rect 52980 64368 53044 64432
rect 53060 64368 53124 64432
rect 53140 64368 53204 64432
rect 53220 64368 53284 64432
rect 58740 64368 58804 64432
rect 58820 64368 58884 64432
rect 58900 64368 58964 64432
rect 58980 64368 59044 64432
rect 59060 64428 59124 64432
rect 59060 64372 59104 64428
rect 59104 64372 59124 64428
rect 59060 64368 59124 64372
rect 59140 64368 59204 64432
rect 59220 64368 59284 64432
rect 64740 64368 64804 64432
rect 64820 64368 64884 64432
rect 64900 64368 64964 64432
rect 64980 64368 65044 64432
rect 65060 64368 65124 64432
rect 65140 64368 65204 64432
rect 65220 64368 65284 64432
rect 70740 64368 70804 64432
rect 70820 64368 70884 64432
rect 70900 64368 70964 64432
rect 70980 64368 71044 64432
rect 71060 64368 71124 64432
rect 71140 64368 71204 64432
rect 71220 64368 71284 64432
rect 4740 64288 4804 64352
rect 4820 64288 4884 64352
rect 4900 64288 4964 64352
rect 4980 64288 5044 64352
rect 5060 64288 5124 64352
rect 5140 64288 5204 64352
rect 5220 64288 5284 64352
rect 10740 64288 10804 64352
rect 10820 64288 10884 64352
rect 10900 64288 10964 64352
rect 10980 64288 11044 64352
rect 11060 64288 11124 64352
rect 11140 64288 11204 64352
rect 11220 64288 11284 64352
rect 16740 64288 16804 64352
rect 16820 64288 16884 64352
rect 16900 64288 16964 64352
rect 16980 64288 17044 64352
rect 17060 64348 17124 64352
rect 17140 64348 17204 64352
rect 17060 64292 17100 64348
rect 17100 64292 17124 64348
rect 17140 64292 17156 64348
rect 17156 64292 17204 64348
rect 17060 64288 17124 64292
rect 17140 64288 17204 64292
rect 17220 64288 17284 64352
rect 22740 64288 22804 64352
rect 22820 64348 22884 64352
rect 22900 64348 22964 64352
rect 22820 64292 22880 64348
rect 22880 64292 22884 64348
rect 22900 64292 22936 64348
rect 22936 64292 22964 64348
rect 22820 64288 22884 64292
rect 22900 64288 22964 64292
rect 22980 64288 23044 64352
rect 23060 64288 23124 64352
rect 23140 64288 23204 64352
rect 23220 64288 23284 64352
rect 28740 64288 28804 64352
rect 28820 64288 28884 64352
rect 28900 64288 28964 64352
rect 28980 64288 29044 64352
rect 29060 64288 29124 64352
rect 29140 64288 29204 64352
rect 29220 64288 29284 64352
rect 34740 64288 34804 64352
rect 34820 64288 34884 64352
rect 34900 64288 34964 64352
rect 34980 64288 35044 64352
rect 35060 64288 35124 64352
rect 35140 64288 35204 64352
rect 35220 64288 35284 64352
rect 40740 64288 40804 64352
rect 40820 64288 40884 64352
rect 40900 64288 40964 64352
rect 40980 64288 41044 64352
rect 41060 64288 41124 64352
rect 41140 64288 41204 64352
rect 41220 64288 41284 64352
rect 46740 64288 46804 64352
rect 46820 64288 46884 64352
rect 46900 64288 46964 64352
rect 46980 64288 47044 64352
rect 47060 64288 47124 64352
rect 47140 64288 47204 64352
rect 47220 64288 47284 64352
rect 52740 64288 52804 64352
rect 52820 64288 52884 64352
rect 52900 64288 52964 64352
rect 52980 64288 53044 64352
rect 53060 64288 53124 64352
rect 53140 64288 53204 64352
rect 53220 64288 53284 64352
rect 58740 64288 58804 64352
rect 58820 64288 58884 64352
rect 58900 64288 58964 64352
rect 58980 64288 59044 64352
rect 59060 64348 59124 64352
rect 59060 64292 59104 64348
rect 59104 64292 59124 64348
rect 59060 64288 59124 64292
rect 59140 64288 59204 64352
rect 59220 64288 59284 64352
rect 64740 64288 64804 64352
rect 64820 64288 64884 64352
rect 64900 64288 64964 64352
rect 64980 64288 65044 64352
rect 65060 64288 65124 64352
rect 65140 64288 65204 64352
rect 65220 64288 65284 64352
rect 70740 64288 70804 64352
rect 70820 64288 70884 64352
rect 70900 64288 70964 64352
rect 70980 64288 71044 64352
rect 71060 64288 71124 64352
rect 71140 64288 71204 64352
rect 71220 64288 71284 64352
rect 1740 62176 1804 62240
rect 1820 62176 1884 62240
rect 1900 62176 1964 62240
rect 1980 62176 2044 62240
rect 2060 62176 2124 62240
rect 2140 62236 2204 62240
rect 2220 62236 2284 62240
rect 2140 62180 2184 62236
rect 2184 62180 2204 62236
rect 2220 62180 2240 62236
rect 2240 62180 2264 62236
rect 2264 62180 2284 62236
rect 2140 62176 2204 62180
rect 2220 62176 2284 62180
rect 7740 62176 7804 62240
rect 7820 62176 7884 62240
rect 7900 62176 7964 62240
rect 7980 62176 8044 62240
rect 8060 62176 8124 62240
rect 8140 62176 8204 62240
rect 8220 62236 8284 62240
rect 8220 62180 8283 62236
rect 8283 62180 8284 62236
rect 8220 62176 8284 62180
rect 13740 62176 13804 62240
rect 13820 62176 13884 62240
rect 13900 62176 13964 62240
rect 13980 62176 14044 62240
rect 14060 62236 14124 62240
rect 14060 62180 14063 62236
rect 14063 62180 14119 62236
rect 14119 62180 14124 62236
rect 14060 62176 14124 62180
rect 14140 62176 14204 62240
rect 14220 62176 14284 62240
rect 19740 62176 19804 62240
rect 19820 62236 19884 62240
rect 19820 62180 19843 62236
rect 19843 62180 19884 62236
rect 19820 62176 19884 62180
rect 19900 62176 19964 62240
rect 19980 62176 20044 62240
rect 20060 62176 20124 62240
rect 20140 62176 20204 62240
rect 20220 62176 20284 62240
rect 25740 62176 25804 62240
rect 25820 62176 25884 62240
rect 25900 62176 25964 62240
rect 25980 62176 26044 62240
rect 26060 62176 26124 62240
rect 26140 62176 26204 62240
rect 26220 62176 26284 62240
rect 31740 62176 31804 62240
rect 31820 62176 31884 62240
rect 31900 62176 31964 62240
rect 31980 62176 32044 62240
rect 32060 62176 32124 62240
rect 32140 62176 32204 62240
rect 32220 62176 32284 62240
rect 37740 62176 37804 62240
rect 37820 62176 37884 62240
rect 37900 62176 37964 62240
rect 37980 62176 38044 62240
rect 38060 62176 38124 62240
rect 38140 62176 38204 62240
rect 38220 62176 38284 62240
rect 43740 62176 43804 62240
rect 43820 62176 43884 62240
rect 43900 62176 43964 62240
rect 43980 62176 44044 62240
rect 44060 62176 44124 62240
rect 44140 62176 44204 62240
rect 44220 62176 44284 62240
rect 49740 62236 49804 62240
rect 49740 62180 49742 62236
rect 49742 62180 49798 62236
rect 49798 62180 49804 62236
rect 49740 62176 49804 62180
rect 49820 62176 49884 62240
rect 49900 62176 49964 62240
rect 49980 62176 50044 62240
rect 50060 62176 50124 62240
rect 50140 62176 50204 62240
rect 50220 62176 50284 62240
rect 55740 62176 55804 62240
rect 55820 62176 55884 62240
rect 55900 62176 55964 62240
rect 55980 62176 56044 62240
rect 56060 62176 56124 62240
rect 56140 62176 56204 62240
rect 56220 62176 56284 62240
rect 61740 62176 61804 62240
rect 61820 62176 61884 62240
rect 61900 62176 61964 62240
rect 61980 62176 62044 62240
rect 62060 62176 62124 62240
rect 62140 62176 62204 62240
rect 62220 62176 62284 62240
rect 67740 62176 67804 62240
rect 67820 62176 67884 62240
rect 67900 62176 67964 62240
rect 67980 62176 68044 62240
rect 68060 62176 68124 62240
rect 68140 62176 68204 62240
rect 68220 62176 68284 62240
rect 73740 62176 73804 62240
rect 73820 62176 73884 62240
rect 73900 62176 73964 62240
rect 73980 62176 74044 62240
rect 74060 62176 74124 62240
rect 74140 62176 74204 62240
rect 74220 62176 74284 62240
rect 1740 62096 1804 62160
rect 1820 62096 1884 62160
rect 1900 62096 1964 62160
rect 1980 62096 2044 62160
rect 2060 62096 2124 62160
rect 2140 62156 2204 62160
rect 2220 62156 2284 62160
rect 2140 62100 2184 62156
rect 2184 62100 2204 62156
rect 2220 62100 2240 62156
rect 2240 62100 2264 62156
rect 2264 62100 2284 62156
rect 2140 62096 2204 62100
rect 2220 62096 2284 62100
rect 7740 62096 7804 62160
rect 7820 62096 7884 62160
rect 7900 62096 7964 62160
rect 7980 62096 8044 62160
rect 8060 62096 8124 62160
rect 8140 62096 8204 62160
rect 8220 62156 8284 62160
rect 8220 62100 8283 62156
rect 8283 62100 8284 62156
rect 8220 62096 8284 62100
rect 13740 62096 13804 62160
rect 13820 62096 13884 62160
rect 13900 62096 13964 62160
rect 13980 62096 14044 62160
rect 14060 62156 14124 62160
rect 14060 62100 14063 62156
rect 14063 62100 14119 62156
rect 14119 62100 14124 62156
rect 14060 62096 14124 62100
rect 14140 62096 14204 62160
rect 14220 62096 14284 62160
rect 19740 62096 19804 62160
rect 19820 62156 19884 62160
rect 19820 62100 19843 62156
rect 19843 62100 19884 62156
rect 19820 62096 19884 62100
rect 19900 62096 19964 62160
rect 19980 62096 20044 62160
rect 20060 62096 20124 62160
rect 20140 62096 20204 62160
rect 20220 62096 20284 62160
rect 25740 62096 25804 62160
rect 25820 62096 25884 62160
rect 25900 62096 25964 62160
rect 25980 62096 26044 62160
rect 26060 62096 26124 62160
rect 26140 62096 26204 62160
rect 26220 62096 26284 62160
rect 31740 62096 31804 62160
rect 31820 62096 31884 62160
rect 31900 62096 31964 62160
rect 31980 62096 32044 62160
rect 32060 62096 32124 62160
rect 32140 62096 32204 62160
rect 32220 62096 32284 62160
rect 37740 62096 37804 62160
rect 37820 62096 37884 62160
rect 37900 62096 37964 62160
rect 37980 62096 38044 62160
rect 38060 62096 38124 62160
rect 38140 62096 38204 62160
rect 38220 62096 38284 62160
rect 43740 62096 43804 62160
rect 43820 62096 43884 62160
rect 43900 62096 43964 62160
rect 43980 62096 44044 62160
rect 44060 62096 44124 62160
rect 44140 62096 44204 62160
rect 44220 62096 44284 62160
rect 49740 62156 49804 62160
rect 49740 62100 49742 62156
rect 49742 62100 49798 62156
rect 49798 62100 49804 62156
rect 49740 62096 49804 62100
rect 49820 62096 49884 62160
rect 49900 62096 49964 62160
rect 49980 62096 50044 62160
rect 50060 62096 50124 62160
rect 50140 62096 50204 62160
rect 50220 62096 50284 62160
rect 55740 62096 55804 62160
rect 55820 62096 55884 62160
rect 55900 62096 55964 62160
rect 55980 62096 56044 62160
rect 56060 62096 56124 62160
rect 56140 62096 56204 62160
rect 56220 62096 56284 62160
rect 61740 62096 61804 62160
rect 61820 62096 61884 62160
rect 61900 62096 61964 62160
rect 61980 62096 62044 62160
rect 62060 62096 62124 62160
rect 62140 62096 62204 62160
rect 62220 62096 62284 62160
rect 67740 62096 67804 62160
rect 67820 62096 67884 62160
rect 67900 62096 67964 62160
rect 67980 62096 68044 62160
rect 68060 62096 68124 62160
rect 68140 62096 68204 62160
rect 68220 62096 68284 62160
rect 73740 62096 73804 62160
rect 73820 62096 73884 62160
rect 73900 62096 73964 62160
rect 73980 62096 74044 62160
rect 74060 62096 74124 62160
rect 74140 62096 74204 62160
rect 74220 62096 74284 62160
rect 1740 62016 1804 62080
rect 1820 62016 1884 62080
rect 1900 62016 1964 62080
rect 1980 62016 2044 62080
rect 2060 62016 2124 62080
rect 2140 62076 2204 62080
rect 2220 62076 2284 62080
rect 2140 62020 2184 62076
rect 2184 62020 2204 62076
rect 2220 62020 2240 62076
rect 2240 62020 2264 62076
rect 2264 62020 2284 62076
rect 2140 62016 2204 62020
rect 2220 62016 2284 62020
rect 7740 62016 7804 62080
rect 7820 62016 7884 62080
rect 7900 62016 7964 62080
rect 7980 62016 8044 62080
rect 8060 62016 8124 62080
rect 8140 62016 8204 62080
rect 8220 62076 8284 62080
rect 8220 62020 8283 62076
rect 8283 62020 8284 62076
rect 8220 62016 8284 62020
rect 13740 62016 13804 62080
rect 13820 62016 13884 62080
rect 13900 62016 13964 62080
rect 13980 62016 14044 62080
rect 14060 62076 14124 62080
rect 14060 62020 14063 62076
rect 14063 62020 14119 62076
rect 14119 62020 14124 62076
rect 14060 62016 14124 62020
rect 14140 62016 14204 62080
rect 14220 62016 14284 62080
rect 19740 62016 19804 62080
rect 19820 62076 19884 62080
rect 19820 62020 19843 62076
rect 19843 62020 19884 62076
rect 19820 62016 19884 62020
rect 19900 62016 19964 62080
rect 19980 62016 20044 62080
rect 20060 62016 20124 62080
rect 20140 62016 20204 62080
rect 20220 62016 20284 62080
rect 25740 62016 25804 62080
rect 25820 62016 25884 62080
rect 25900 62016 25964 62080
rect 25980 62016 26044 62080
rect 26060 62016 26124 62080
rect 26140 62016 26204 62080
rect 26220 62016 26284 62080
rect 31740 62016 31804 62080
rect 31820 62016 31884 62080
rect 31900 62016 31964 62080
rect 31980 62016 32044 62080
rect 32060 62016 32124 62080
rect 32140 62016 32204 62080
rect 32220 62016 32284 62080
rect 37740 62016 37804 62080
rect 37820 62016 37884 62080
rect 37900 62016 37964 62080
rect 37980 62016 38044 62080
rect 38060 62016 38124 62080
rect 38140 62016 38204 62080
rect 38220 62016 38284 62080
rect 43740 62016 43804 62080
rect 43820 62016 43884 62080
rect 43900 62016 43964 62080
rect 43980 62016 44044 62080
rect 44060 62016 44124 62080
rect 44140 62016 44204 62080
rect 44220 62016 44284 62080
rect 49740 62076 49804 62080
rect 49740 62020 49742 62076
rect 49742 62020 49798 62076
rect 49798 62020 49804 62076
rect 49740 62016 49804 62020
rect 49820 62016 49884 62080
rect 49900 62016 49964 62080
rect 49980 62016 50044 62080
rect 50060 62016 50124 62080
rect 50140 62016 50204 62080
rect 50220 62016 50284 62080
rect 55740 62016 55804 62080
rect 55820 62016 55884 62080
rect 55900 62016 55964 62080
rect 55980 62016 56044 62080
rect 56060 62016 56124 62080
rect 56140 62016 56204 62080
rect 56220 62016 56284 62080
rect 61740 62016 61804 62080
rect 61820 62016 61884 62080
rect 61900 62016 61964 62080
rect 61980 62016 62044 62080
rect 62060 62016 62124 62080
rect 62140 62016 62204 62080
rect 62220 62016 62284 62080
rect 67740 62016 67804 62080
rect 67820 62016 67884 62080
rect 67900 62016 67964 62080
rect 67980 62016 68044 62080
rect 68060 62016 68124 62080
rect 68140 62016 68204 62080
rect 68220 62016 68284 62080
rect 73740 62016 73804 62080
rect 73820 62016 73884 62080
rect 73900 62016 73964 62080
rect 73980 62016 74044 62080
rect 74060 62016 74124 62080
rect 74140 62016 74204 62080
rect 74220 62016 74284 62080
rect 1740 61936 1804 62000
rect 1820 61936 1884 62000
rect 1900 61936 1964 62000
rect 1980 61936 2044 62000
rect 2060 61936 2124 62000
rect 2140 61996 2204 62000
rect 2220 61996 2284 62000
rect 2140 61940 2184 61996
rect 2184 61940 2204 61996
rect 2220 61940 2240 61996
rect 2240 61940 2264 61996
rect 2264 61940 2284 61996
rect 2140 61936 2204 61940
rect 2220 61936 2284 61940
rect 7740 61936 7804 62000
rect 7820 61936 7884 62000
rect 7900 61936 7964 62000
rect 7980 61936 8044 62000
rect 8060 61936 8124 62000
rect 8140 61936 8204 62000
rect 8220 61996 8284 62000
rect 8220 61940 8283 61996
rect 8283 61940 8284 61996
rect 8220 61936 8284 61940
rect 13740 61936 13804 62000
rect 13820 61936 13884 62000
rect 13900 61936 13964 62000
rect 13980 61936 14044 62000
rect 14060 61996 14124 62000
rect 14060 61940 14063 61996
rect 14063 61940 14119 61996
rect 14119 61940 14124 61996
rect 14060 61936 14124 61940
rect 14140 61936 14204 62000
rect 14220 61936 14284 62000
rect 19740 61936 19804 62000
rect 19820 61996 19884 62000
rect 19820 61940 19843 61996
rect 19843 61940 19884 61996
rect 19820 61936 19884 61940
rect 19900 61936 19964 62000
rect 19980 61936 20044 62000
rect 20060 61936 20124 62000
rect 20140 61936 20204 62000
rect 20220 61936 20284 62000
rect 25740 61936 25804 62000
rect 25820 61936 25884 62000
rect 25900 61936 25964 62000
rect 25980 61936 26044 62000
rect 26060 61936 26124 62000
rect 26140 61936 26204 62000
rect 26220 61936 26284 62000
rect 31740 61936 31804 62000
rect 31820 61936 31884 62000
rect 31900 61936 31964 62000
rect 31980 61936 32044 62000
rect 32060 61936 32124 62000
rect 32140 61936 32204 62000
rect 32220 61936 32284 62000
rect 37740 61936 37804 62000
rect 37820 61936 37884 62000
rect 37900 61936 37964 62000
rect 37980 61936 38044 62000
rect 38060 61936 38124 62000
rect 38140 61936 38204 62000
rect 38220 61936 38284 62000
rect 43740 61936 43804 62000
rect 43820 61936 43884 62000
rect 43900 61936 43964 62000
rect 43980 61936 44044 62000
rect 44060 61936 44124 62000
rect 44140 61936 44204 62000
rect 44220 61936 44284 62000
rect 49740 61996 49804 62000
rect 49740 61940 49742 61996
rect 49742 61940 49798 61996
rect 49798 61940 49804 61996
rect 49740 61936 49804 61940
rect 49820 61936 49884 62000
rect 49900 61936 49964 62000
rect 49980 61936 50044 62000
rect 50060 61936 50124 62000
rect 50140 61936 50204 62000
rect 50220 61936 50284 62000
rect 55740 61936 55804 62000
rect 55820 61936 55884 62000
rect 55900 61936 55964 62000
rect 55980 61936 56044 62000
rect 56060 61936 56124 62000
rect 56140 61936 56204 62000
rect 56220 61936 56284 62000
rect 61740 61936 61804 62000
rect 61820 61936 61884 62000
rect 61900 61936 61964 62000
rect 61980 61936 62044 62000
rect 62060 61936 62124 62000
rect 62140 61936 62204 62000
rect 62220 61936 62284 62000
rect 67740 61936 67804 62000
rect 67820 61936 67884 62000
rect 67900 61936 67964 62000
rect 67980 61936 68044 62000
rect 68060 61936 68124 62000
rect 68140 61936 68204 62000
rect 68220 61936 68284 62000
rect 73740 61936 73804 62000
rect 73820 61936 73884 62000
rect 73900 61936 73964 62000
rect 73980 61936 74044 62000
rect 74060 61936 74124 62000
rect 74140 61936 74204 62000
rect 74220 61936 74284 62000
rect 4740 54528 4804 54592
rect 4820 54528 4884 54592
rect 4900 54528 4964 54592
rect 4980 54528 5044 54592
rect 5060 54528 5124 54592
rect 5140 54528 5204 54592
rect 5220 54528 5284 54592
rect 10740 54528 10804 54592
rect 10820 54528 10884 54592
rect 10900 54528 10964 54592
rect 10980 54528 11044 54592
rect 11060 54528 11124 54592
rect 11140 54528 11204 54592
rect 11220 54528 11284 54592
rect 16740 54528 16804 54592
rect 16820 54528 16884 54592
rect 16900 54528 16964 54592
rect 16980 54528 17044 54592
rect 17060 54588 17124 54592
rect 17140 54588 17204 54592
rect 17060 54532 17100 54588
rect 17100 54532 17124 54588
rect 17140 54532 17156 54588
rect 17156 54532 17204 54588
rect 17060 54528 17124 54532
rect 17140 54528 17204 54532
rect 17220 54528 17284 54592
rect 22740 54528 22804 54592
rect 22820 54588 22884 54592
rect 22900 54588 22964 54592
rect 22820 54532 22880 54588
rect 22880 54532 22884 54588
rect 22900 54532 22936 54588
rect 22936 54532 22964 54588
rect 22820 54528 22884 54532
rect 22900 54528 22964 54532
rect 22980 54528 23044 54592
rect 23060 54528 23124 54592
rect 23140 54528 23204 54592
rect 23220 54528 23284 54592
rect 28740 54528 28804 54592
rect 28820 54528 28884 54592
rect 28900 54528 28964 54592
rect 28980 54528 29044 54592
rect 29060 54528 29124 54592
rect 29140 54528 29204 54592
rect 29220 54528 29284 54592
rect 34740 54528 34804 54592
rect 34820 54528 34884 54592
rect 34900 54528 34964 54592
rect 34980 54528 35044 54592
rect 35060 54528 35124 54592
rect 35140 54528 35204 54592
rect 35220 54528 35284 54592
rect 40740 54528 40804 54592
rect 40820 54528 40884 54592
rect 40900 54528 40964 54592
rect 40980 54528 41044 54592
rect 41060 54528 41124 54592
rect 41140 54528 41204 54592
rect 41220 54528 41284 54592
rect 46740 54528 46804 54592
rect 46820 54528 46884 54592
rect 46900 54528 46964 54592
rect 46980 54528 47044 54592
rect 47060 54528 47124 54592
rect 47140 54528 47204 54592
rect 47220 54528 47284 54592
rect 52740 54528 52804 54592
rect 52820 54528 52884 54592
rect 52900 54528 52964 54592
rect 52980 54528 53044 54592
rect 53060 54528 53124 54592
rect 53140 54528 53204 54592
rect 53220 54528 53284 54592
rect 58740 54528 58804 54592
rect 58820 54528 58884 54592
rect 58900 54528 58964 54592
rect 58980 54528 59044 54592
rect 59060 54588 59124 54592
rect 59060 54532 59104 54588
rect 59104 54532 59124 54588
rect 59060 54528 59124 54532
rect 59140 54528 59204 54592
rect 59220 54528 59284 54592
rect 64740 54528 64804 54592
rect 64820 54528 64884 54592
rect 64900 54528 64964 54592
rect 64980 54528 65044 54592
rect 65060 54528 65124 54592
rect 65140 54528 65204 54592
rect 65220 54528 65284 54592
rect 70740 54528 70804 54592
rect 70820 54528 70884 54592
rect 70900 54528 70964 54592
rect 70980 54528 71044 54592
rect 71060 54528 71124 54592
rect 71140 54528 71204 54592
rect 71220 54528 71284 54592
rect 4740 54448 4804 54512
rect 4820 54448 4884 54512
rect 4900 54448 4964 54512
rect 4980 54448 5044 54512
rect 5060 54448 5124 54512
rect 5140 54448 5204 54512
rect 5220 54448 5284 54512
rect 10740 54448 10804 54512
rect 10820 54448 10884 54512
rect 10900 54448 10964 54512
rect 10980 54448 11044 54512
rect 11060 54448 11124 54512
rect 11140 54448 11204 54512
rect 11220 54448 11284 54512
rect 16740 54448 16804 54512
rect 16820 54448 16884 54512
rect 16900 54448 16964 54512
rect 16980 54448 17044 54512
rect 17060 54508 17124 54512
rect 17140 54508 17204 54512
rect 17060 54452 17100 54508
rect 17100 54452 17124 54508
rect 17140 54452 17156 54508
rect 17156 54452 17204 54508
rect 17060 54448 17124 54452
rect 17140 54448 17204 54452
rect 17220 54448 17284 54512
rect 22740 54448 22804 54512
rect 22820 54508 22884 54512
rect 22900 54508 22964 54512
rect 22820 54452 22880 54508
rect 22880 54452 22884 54508
rect 22900 54452 22936 54508
rect 22936 54452 22964 54508
rect 22820 54448 22884 54452
rect 22900 54448 22964 54452
rect 22980 54448 23044 54512
rect 23060 54448 23124 54512
rect 23140 54448 23204 54512
rect 23220 54448 23284 54512
rect 28740 54448 28804 54512
rect 28820 54448 28884 54512
rect 28900 54448 28964 54512
rect 28980 54448 29044 54512
rect 29060 54448 29124 54512
rect 29140 54448 29204 54512
rect 29220 54448 29284 54512
rect 34740 54448 34804 54512
rect 34820 54448 34884 54512
rect 34900 54448 34964 54512
rect 34980 54448 35044 54512
rect 35060 54448 35124 54512
rect 35140 54448 35204 54512
rect 35220 54448 35284 54512
rect 40740 54448 40804 54512
rect 40820 54448 40884 54512
rect 40900 54448 40964 54512
rect 40980 54448 41044 54512
rect 41060 54448 41124 54512
rect 41140 54448 41204 54512
rect 41220 54448 41284 54512
rect 46740 54448 46804 54512
rect 46820 54448 46884 54512
rect 46900 54448 46964 54512
rect 46980 54448 47044 54512
rect 47060 54448 47124 54512
rect 47140 54448 47204 54512
rect 47220 54448 47284 54512
rect 52740 54448 52804 54512
rect 52820 54448 52884 54512
rect 52900 54448 52964 54512
rect 52980 54448 53044 54512
rect 53060 54448 53124 54512
rect 53140 54448 53204 54512
rect 53220 54448 53284 54512
rect 58740 54448 58804 54512
rect 58820 54448 58884 54512
rect 58900 54448 58964 54512
rect 58980 54448 59044 54512
rect 59060 54508 59124 54512
rect 59060 54452 59104 54508
rect 59104 54452 59124 54508
rect 59060 54448 59124 54452
rect 59140 54448 59204 54512
rect 59220 54448 59284 54512
rect 64740 54448 64804 54512
rect 64820 54448 64884 54512
rect 64900 54448 64964 54512
rect 64980 54448 65044 54512
rect 65060 54448 65124 54512
rect 65140 54448 65204 54512
rect 65220 54448 65284 54512
rect 70740 54448 70804 54512
rect 70820 54448 70884 54512
rect 70900 54448 70964 54512
rect 70980 54448 71044 54512
rect 71060 54448 71124 54512
rect 71140 54448 71204 54512
rect 71220 54448 71284 54512
rect 4740 54368 4804 54432
rect 4820 54368 4884 54432
rect 4900 54368 4964 54432
rect 4980 54368 5044 54432
rect 5060 54368 5124 54432
rect 5140 54368 5204 54432
rect 5220 54368 5284 54432
rect 10740 54368 10804 54432
rect 10820 54368 10884 54432
rect 10900 54368 10964 54432
rect 10980 54368 11044 54432
rect 11060 54368 11124 54432
rect 11140 54368 11204 54432
rect 11220 54368 11284 54432
rect 16740 54368 16804 54432
rect 16820 54368 16884 54432
rect 16900 54368 16964 54432
rect 16980 54368 17044 54432
rect 17060 54428 17124 54432
rect 17140 54428 17204 54432
rect 17060 54372 17100 54428
rect 17100 54372 17124 54428
rect 17140 54372 17156 54428
rect 17156 54372 17204 54428
rect 17060 54368 17124 54372
rect 17140 54368 17204 54372
rect 17220 54368 17284 54432
rect 22740 54368 22804 54432
rect 22820 54428 22884 54432
rect 22900 54428 22964 54432
rect 22820 54372 22880 54428
rect 22880 54372 22884 54428
rect 22900 54372 22936 54428
rect 22936 54372 22964 54428
rect 22820 54368 22884 54372
rect 22900 54368 22964 54372
rect 22980 54368 23044 54432
rect 23060 54368 23124 54432
rect 23140 54368 23204 54432
rect 23220 54368 23284 54432
rect 28740 54368 28804 54432
rect 28820 54368 28884 54432
rect 28900 54368 28964 54432
rect 28980 54368 29044 54432
rect 29060 54368 29124 54432
rect 29140 54368 29204 54432
rect 29220 54368 29284 54432
rect 34740 54368 34804 54432
rect 34820 54368 34884 54432
rect 34900 54368 34964 54432
rect 34980 54368 35044 54432
rect 35060 54368 35124 54432
rect 35140 54368 35204 54432
rect 35220 54368 35284 54432
rect 40740 54368 40804 54432
rect 40820 54368 40884 54432
rect 40900 54368 40964 54432
rect 40980 54368 41044 54432
rect 41060 54368 41124 54432
rect 41140 54368 41204 54432
rect 41220 54368 41284 54432
rect 46740 54368 46804 54432
rect 46820 54368 46884 54432
rect 46900 54368 46964 54432
rect 46980 54368 47044 54432
rect 47060 54368 47124 54432
rect 47140 54368 47204 54432
rect 47220 54368 47284 54432
rect 52740 54368 52804 54432
rect 52820 54368 52884 54432
rect 52900 54368 52964 54432
rect 52980 54368 53044 54432
rect 53060 54368 53124 54432
rect 53140 54368 53204 54432
rect 53220 54368 53284 54432
rect 58740 54368 58804 54432
rect 58820 54368 58884 54432
rect 58900 54368 58964 54432
rect 58980 54368 59044 54432
rect 59060 54428 59124 54432
rect 59060 54372 59104 54428
rect 59104 54372 59124 54428
rect 59060 54368 59124 54372
rect 59140 54368 59204 54432
rect 59220 54368 59284 54432
rect 64740 54368 64804 54432
rect 64820 54368 64884 54432
rect 64900 54368 64964 54432
rect 64980 54368 65044 54432
rect 65060 54368 65124 54432
rect 65140 54368 65204 54432
rect 65220 54368 65284 54432
rect 70740 54368 70804 54432
rect 70820 54368 70884 54432
rect 70900 54368 70964 54432
rect 70980 54368 71044 54432
rect 71060 54368 71124 54432
rect 71140 54368 71204 54432
rect 71220 54368 71284 54432
rect 4740 54288 4804 54352
rect 4820 54288 4884 54352
rect 4900 54288 4964 54352
rect 4980 54288 5044 54352
rect 5060 54288 5124 54352
rect 5140 54288 5204 54352
rect 5220 54288 5284 54352
rect 10740 54288 10804 54352
rect 10820 54288 10884 54352
rect 10900 54288 10964 54352
rect 10980 54288 11044 54352
rect 11060 54288 11124 54352
rect 11140 54288 11204 54352
rect 11220 54288 11284 54352
rect 16740 54288 16804 54352
rect 16820 54288 16884 54352
rect 16900 54288 16964 54352
rect 16980 54288 17044 54352
rect 17060 54348 17124 54352
rect 17140 54348 17204 54352
rect 17060 54292 17100 54348
rect 17100 54292 17124 54348
rect 17140 54292 17156 54348
rect 17156 54292 17204 54348
rect 17060 54288 17124 54292
rect 17140 54288 17204 54292
rect 17220 54288 17284 54352
rect 22740 54288 22804 54352
rect 22820 54348 22884 54352
rect 22900 54348 22964 54352
rect 22820 54292 22880 54348
rect 22880 54292 22884 54348
rect 22900 54292 22936 54348
rect 22936 54292 22964 54348
rect 22820 54288 22884 54292
rect 22900 54288 22964 54292
rect 22980 54288 23044 54352
rect 23060 54288 23124 54352
rect 23140 54288 23204 54352
rect 23220 54288 23284 54352
rect 28740 54288 28804 54352
rect 28820 54288 28884 54352
rect 28900 54288 28964 54352
rect 28980 54288 29044 54352
rect 29060 54288 29124 54352
rect 29140 54288 29204 54352
rect 29220 54288 29284 54352
rect 34740 54288 34804 54352
rect 34820 54288 34884 54352
rect 34900 54288 34964 54352
rect 34980 54288 35044 54352
rect 35060 54288 35124 54352
rect 35140 54288 35204 54352
rect 35220 54288 35284 54352
rect 40740 54288 40804 54352
rect 40820 54288 40884 54352
rect 40900 54288 40964 54352
rect 40980 54288 41044 54352
rect 41060 54288 41124 54352
rect 41140 54288 41204 54352
rect 41220 54288 41284 54352
rect 46740 54288 46804 54352
rect 46820 54288 46884 54352
rect 46900 54288 46964 54352
rect 46980 54288 47044 54352
rect 47060 54288 47124 54352
rect 47140 54288 47204 54352
rect 47220 54288 47284 54352
rect 52740 54288 52804 54352
rect 52820 54288 52884 54352
rect 52900 54288 52964 54352
rect 52980 54288 53044 54352
rect 53060 54288 53124 54352
rect 53140 54288 53204 54352
rect 53220 54288 53284 54352
rect 58740 54288 58804 54352
rect 58820 54288 58884 54352
rect 58900 54288 58964 54352
rect 58980 54288 59044 54352
rect 59060 54348 59124 54352
rect 59060 54292 59104 54348
rect 59104 54292 59124 54348
rect 59060 54288 59124 54292
rect 59140 54288 59204 54352
rect 59220 54288 59284 54352
rect 64740 54288 64804 54352
rect 64820 54288 64884 54352
rect 64900 54288 64964 54352
rect 64980 54288 65044 54352
rect 65060 54288 65124 54352
rect 65140 54288 65204 54352
rect 65220 54288 65284 54352
rect 70740 54288 70804 54352
rect 70820 54288 70884 54352
rect 70900 54288 70964 54352
rect 70980 54288 71044 54352
rect 71060 54288 71124 54352
rect 71140 54288 71204 54352
rect 71220 54288 71284 54352
rect 64092 52532 64156 52596
rect 1740 52176 1804 52240
rect 1820 52176 1884 52240
rect 1900 52176 1964 52240
rect 1980 52176 2044 52240
rect 2060 52176 2124 52240
rect 2140 52236 2204 52240
rect 2220 52236 2284 52240
rect 2140 52180 2184 52236
rect 2184 52180 2204 52236
rect 2220 52180 2240 52236
rect 2240 52180 2264 52236
rect 2264 52180 2284 52236
rect 2140 52176 2204 52180
rect 2220 52176 2284 52180
rect 7740 52176 7804 52240
rect 7820 52176 7884 52240
rect 7900 52176 7964 52240
rect 7980 52176 8044 52240
rect 8060 52176 8124 52240
rect 8140 52176 8204 52240
rect 8220 52236 8284 52240
rect 8220 52180 8283 52236
rect 8283 52180 8284 52236
rect 8220 52176 8284 52180
rect 13740 52176 13804 52240
rect 13820 52176 13884 52240
rect 13900 52176 13964 52240
rect 13980 52176 14044 52240
rect 14060 52236 14124 52240
rect 14060 52180 14063 52236
rect 14063 52180 14119 52236
rect 14119 52180 14124 52236
rect 14060 52176 14124 52180
rect 14140 52176 14204 52240
rect 14220 52176 14284 52240
rect 19740 52176 19804 52240
rect 19820 52236 19884 52240
rect 19820 52180 19843 52236
rect 19843 52180 19884 52236
rect 19820 52176 19884 52180
rect 19900 52176 19964 52240
rect 19980 52176 20044 52240
rect 20060 52176 20124 52240
rect 20140 52176 20204 52240
rect 20220 52176 20284 52240
rect 25740 52176 25804 52240
rect 25820 52176 25884 52240
rect 25900 52176 25964 52240
rect 25980 52176 26044 52240
rect 26060 52176 26124 52240
rect 26140 52176 26204 52240
rect 26220 52176 26284 52240
rect 31740 52176 31804 52240
rect 31820 52176 31884 52240
rect 31900 52176 31964 52240
rect 31980 52176 32044 52240
rect 32060 52176 32124 52240
rect 32140 52176 32204 52240
rect 32220 52176 32284 52240
rect 37740 52176 37804 52240
rect 37820 52176 37884 52240
rect 37900 52176 37964 52240
rect 37980 52176 38044 52240
rect 38060 52176 38124 52240
rect 38140 52176 38204 52240
rect 38220 52176 38284 52240
rect 43740 52176 43804 52240
rect 43820 52176 43884 52240
rect 43900 52176 43964 52240
rect 43980 52176 44044 52240
rect 44060 52176 44124 52240
rect 44140 52176 44204 52240
rect 44220 52176 44284 52240
rect 49740 52236 49804 52240
rect 49740 52180 49742 52236
rect 49742 52180 49798 52236
rect 49798 52180 49804 52236
rect 49740 52176 49804 52180
rect 49820 52176 49884 52240
rect 49900 52176 49964 52240
rect 49980 52176 50044 52240
rect 50060 52176 50124 52240
rect 50140 52176 50204 52240
rect 50220 52176 50284 52240
rect 55740 52176 55804 52240
rect 55820 52176 55884 52240
rect 55900 52176 55964 52240
rect 55980 52176 56044 52240
rect 56060 52176 56124 52240
rect 56140 52176 56204 52240
rect 56220 52176 56284 52240
rect 61740 52176 61804 52240
rect 61820 52176 61884 52240
rect 61900 52176 61964 52240
rect 61980 52176 62044 52240
rect 62060 52176 62124 52240
rect 62140 52176 62204 52240
rect 62220 52176 62284 52240
rect 67740 52176 67804 52240
rect 67820 52176 67884 52240
rect 67900 52176 67964 52240
rect 67980 52176 68044 52240
rect 68060 52176 68124 52240
rect 68140 52176 68204 52240
rect 68220 52176 68284 52240
rect 73740 52176 73804 52240
rect 73820 52176 73884 52240
rect 73900 52176 73964 52240
rect 73980 52176 74044 52240
rect 74060 52176 74124 52240
rect 74140 52176 74204 52240
rect 74220 52176 74284 52240
rect 1740 52096 1804 52160
rect 1820 52096 1884 52160
rect 1900 52096 1964 52160
rect 1980 52096 2044 52160
rect 2060 52096 2124 52160
rect 2140 52156 2204 52160
rect 2220 52156 2284 52160
rect 2140 52100 2184 52156
rect 2184 52100 2204 52156
rect 2220 52100 2240 52156
rect 2240 52100 2264 52156
rect 2264 52100 2284 52156
rect 2140 52096 2204 52100
rect 2220 52096 2284 52100
rect 7740 52096 7804 52160
rect 7820 52096 7884 52160
rect 7900 52096 7964 52160
rect 7980 52096 8044 52160
rect 8060 52096 8124 52160
rect 8140 52096 8204 52160
rect 8220 52156 8284 52160
rect 8220 52100 8283 52156
rect 8283 52100 8284 52156
rect 8220 52096 8284 52100
rect 13740 52096 13804 52160
rect 13820 52096 13884 52160
rect 13900 52096 13964 52160
rect 13980 52096 14044 52160
rect 14060 52156 14124 52160
rect 14060 52100 14063 52156
rect 14063 52100 14119 52156
rect 14119 52100 14124 52156
rect 14060 52096 14124 52100
rect 14140 52096 14204 52160
rect 14220 52096 14284 52160
rect 19740 52096 19804 52160
rect 19820 52156 19884 52160
rect 19820 52100 19843 52156
rect 19843 52100 19884 52156
rect 19820 52096 19884 52100
rect 19900 52096 19964 52160
rect 19980 52096 20044 52160
rect 20060 52096 20124 52160
rect 20140 52096 20204 52160
rect 20220 52096 20284 52160
rect 25740 52096 25804 52160
rect 25820 52096 25884 52160
rect 25900 52096 25964 52160
rect 25980 52096 26044 52160
rect 26060 52096 26124 52160
rect 26140 52096 26204 52160
rect 26220 52096 26284 52160
rect 31740 52096 31804 52160
rect 31820 52096 31884 52160
rect 31900 52096 31964 52160
rect 31980 52096 32044 52160
rect 32060 52096 32124 52160
rect 32140 52096 32204 52160
rect 32220 52096 32284 52160
rect 37740 52096 37804 52160
rect 37820 52096 37884 52160
rect 37900 52096 37964 52160
rect 37980 52096 38044 52160
rect 38060 52096 38124 52160
rect 38140 52096 38204 52160
rect 38220 52096 38284 52160
rect 43740 52096 43804 52160
rect 43820 52096 43884 52160
rect 43900 52096 43964 52160
rect 43980 52096 44044 52160
rect 44060 52096 44124 52160
rect 44140 52096 44204 52160
rect 44220 52096 44284 52160
rect 49740 52156 49804 52160
rect 49740 52100 49742 52156
rect 49742 52100 49798 52156
rect 49798 52100 49804 52156
rect 49740 52096 49804 52100
rect 49820 52096 49884 52160
rect 49900 52096 49964 52160
rect 49980 52096 50044 52160
rect 50060 52096 50124 52160
rect 50140 52096 50204 52160
rect 50220 52096 50284 52160
rect 55740 52096 55804 52160
rect 55820 52096 55884 52160
rect 55900 52096 55964 52160
rect 55980 52096 56044 52160
rect 56060 52096 56124 52160
rect 56140 52096 56204 52160
rect 56220 52096 56284 52160
rect 61740 52096 61804 52160
rect 61820 52096 61884 52160
rect 61900 52096 61964 52160
rect 61980 52096 62044 52160
rect 62060 52096 62124 52160
rect 62140 52096 62204 52160
rect 62220 52096 62284 52160
rect 67740 52096 67804 52160
rect 67820 52096 67884 52160
rect 67900 52096 67964 52160
rect 67980 52096 68044 52160
rect 68060 52096 68124 52160
rect 68140 52096 68204 52160
rect 68220 52096 68284 52160
rect 73740 52096 73804 52160
rect 73820 52096 73884 52160
rect 73900 52096 73964 52160
rect 73980 52096 74044 52160
rect 74060 52096 74124 52160
rect 74140 52096 74204 52160
rect 74220 52096 74284 52160
rect 1740 52016 1804 52080
rect 1820 52016 1884 52080
rect 1900 52016 1964 52080
rect 1980 52016 2044 52080
rect 2060 52016 2124 52080
rect 2140 52076 2204 52080
rect 2220 52076 2284 52080
rect 2140 52020 2184 52076
rect 2184 52020 2204 52076
rect 2220 52020 2240 52076
rect 2240 52020 2264 52076
rect 2264 52020 2284 52076
rect 2140 52016 2204 52020
rect 2220 52016 2284 52020
rect 7740 52016 7804 52080
rect 7820 52016 7884 52080
rect 7900 52016 7964 52080
rect 7980 52016 8044 52080
rect 8060 52016 8124 52080
rect 8140 52016 8204 52080
rect 8220 52076 8284 52080
rect 8220 52020 8283 52076
rect 8283 52020 8284 52076
rect 8220 52016 8284 52020
rect 13740 52016 13804 52080
rect 13820 52016 13884 52080
rect 13900 52016 13964 52080
rect 13980 52016 14044 52080
rect 14060 52076 14124 52080
rect 14060 52020 14063 52076
rect 14063 52020 14119 52076
rect 14119 52020 14124 52076
rect 14060 52016 14124 52020
rect 14140 52016 14204 52080
rect 14220 52016 14284 52080
rect 19740 52016 19804 52080
rect 19820 52076 19884 52080
rect 19820 52020 19843 52076
rect 19843 52020 19884 52076
rect 19820 52016 19884 52020
rect 19900 52016 19964 52080
rect 19980 52016 20044 52080
rect 20060 52016 20124 52080
rect 20140 52016 20204 52080
rect 20220 52016 20284 52080
rect 25740 52016 25804 52080
rect 25820 52016 25884 52080
rect 25900 52016 25964 52080
rect 25980 52016 26044 52080
rect 26060 52016 26124 52080
rect 26140 52016 26204 52080
rect 26220 52016 26284 52080
rect 31740 52016 31804 52080
rect 31820 52016 31884 52080
rect 31900 52016 31964 52080
rect 31980 52016 32044 52080
rect 32060 52016 32124 52080
rect 32140 52016 32204 52080
rect 32220 52016 32284 52080
rect 37740 52016 37804 52080
rect 37820 52016 37884 52080
rect 37900 52016 37964 52080
rect 37980 52016 38044 52080
rect 38060 52016 38124 52080
rect 38140 52016 38204 52080
rect 38220 52016 38284 52080
rect 43740 52016 43804 52080
rect 43820 52016 43884 52080
rect 43900 52016 43964 52080
rect 43980 52016 44044 52080
rect 44060 52016 44124 52080
rect 44140 52016 44204 52080
rect 44220 52016 44284 52080
rect 49740 52076 49804 52080
rect 49740 52020 49742 52076
rect 49742 52020 49798 52076
rect 49798 52020 49804 52076
rect 49740 52016 49804 52020
rect 49820 52016 49884 52080
rect 49900 52016 49964 52080
rect 49980 52016 50044 52080
rect 50060 52016 50124 52080
rect 50140 52016 50204 52080
rect 50220 52016 50284 52080
rect 55740 52016 55804 52080
rect 55820 52016 55884 52080
rect 55900 52016 55964 52080
rect 55980 52016 56044 52080
rect 56060 52016 56124 52080
rect 56140 52016 56204 52080
rect 56220 52016 56284 52080
rect 61740 52016 61804 52080
rect 61820 52016 61884 52080
rect 61900 52016 61964 52080
rect 61980 52016 62044 52080
rect 62060 52016 62124 52080
rect 62140 52016 62204 52080
rect 62220 52016 62284 52080
rect 67740 52016 67804 52080
rect 67820 52016 67884 52080
rect 67900 52016 67964 52080
rect 67980 52016 68044 52080
rect 68060 52016 68124 52080
rect 68140 52016 68204 52080
rect 68220 52016 68284 52080
rect 73740 52016 73804 52080
rect 73820 52016 73884 52080
rect 73900 52016 73964 52080
rect 73980 52016 74044 52080
rect 74060 52016 74124 52080
rect 74140 52016 74204 52080
rect 74220 52016 74284 52080
rect 1740 51936 1804 52000
rect 1820 51936 1884 52000
rect 1900 51936 1964 52000
rect 1980 51936 2044 52000
rect 2060 51936 2124 52000
rect 2140 51996 2204 52000
rect 2220 51996 2284 52000
rect 2140 51940 2184 51996
rect 2184 51940 2204 51996
rect 2220 51940 2240 51996
rect 2240 51940 2264 51996
rect 2264 51940 2284 51996
rect 2140 51936 2204 51940
rect 2220 51936 2284 51940
rect 7740 51936 7804 52000
rect 7820 51936 7884 52000
rect 7900 51936 7964 52000
rect 7980 51936 8044 52000
rect 8060 51936 8124 52000
rect 8140 51936 8204 52000
rect 8220 51996 8284 52000
rect 8220 51940 8283 51996
rect 8283 51940 8284 51996
rect 8220 51936 8284 51940
rect 13740 51936 13804 52000
rect 13820 51936 13884 52000
rect 13900 51936 13964 52000
rect 13980 51936 14044 52000
rect 14060 51996 14124 52000
rect 14060 51940 14063 51996
rect 14063 51940 14119 51996
rect 14119 51940 14124 51996
rect 14060 51936 14124 51940
rect 14140 51936 14204 52000
rect 14220 51936 14284 52000
rect 19740 51936 19804 52000
rect 19820 51996 19884 52000
rect 19820 51940 19843 51996
rect 19843 51940 19884 51996
rect 19820 51936 19884 51940
rect 19900 51936 19964 52000
rect 19980 51936 20044 52000
rect 20060 51936 20124 52000
rect 20140 51936 20204 52000
rect 20220 51936 20284 52000
rect 25740 51936 25804 52000
rect 25820 51936 25884 52000
rect 25900 51936 25964 52000
rect 25980 51936 26044 52000
rect 26060 51936 26124 52000
rect 26140 51936 26204 52000
rect 26220 51936 26284 52000
rect 31740 51936 31804 52000
rect 31820 51936 31884 52000
rect 31900 51936 31964 52000
rect 31980 51936 32044 52000
rect 32060 51936 32124 52000
rect 32140 51936 32204 52000
rect 32220 51936 32284 52000
rect 37740 51936 37804 52000
rect 37820 51936 37884 52000
rect 37900 51936 37964 52000
rect 37980 51936 38044 52000
rect 38060 51936 38124 52000
rect 38140 51936 38204 52000
rect 38220 51936 38284 52000
rect 43740 51936 43804 52000
rect 43820 51936 43884 52000
rect 43900 51936 43964 52000
rect 43980 51936 44044 52000
rect 44060 51936 44124 52000
rect 44140 51936 44204 52000
rect 44220 51936 44284 52000
rect 49740 51996 49804 52000
rect 49740 51940 49742 51996
rect 49742 51940 49798 51996
rect 49798 51940 49804 51996
rect 49740 51936 49804 51940
rect 49820 51936 49884 52000
rect 49900 51936 49964 52000
rect 49980 51936 50044 52000
rect 50060 51936 50124 52000
rect 50140 51936 50204 52000
rect 50220 51936 50284 52000
rect 55740 51936 55804 52000
rect 55820 51936 55884 52000
rect 55900 51936 55964 52000
rect 55980 51936 56044 52000
rect 56060 51936 56124 52000
rect 56140 51936 56204 52000
rect 56220 51936 56284 52000
rect 61740 51936 61804 52000
rect 61820 51936 61884 52000
rect 61900 51936 61964 52000
rect 61980 51936 62044 52000
rect 62060 51936 62124 52000
rect 62140 51936 62204 52000
rect 62220 51936 62284 52000
rect 67740 51936 67804 52000
rect 67820 51936 67884 52000
rect 67900 51936 67964 52000
rect 67980 51936 68044 52000
rect 68060 51936 68124 52000
rect 68140 51936 68204 52000
rect 68220 51936 68284 52000
rect 73740 51936 73804 52000
rect 73820 51936 73884 52000
rect 73900 51936 73964 52000
rect 73980 51936 74044 52000
rect 74060 51936 74124 52000
rect 74140 51936 74204 52000
rect 74220 51936 74284 52000
rect 64276 50220 64340 50284
rect 65564 48044 65628 48108
rect 64460 47696 64524 47700
rect 64460 47640 64474 47696
rect 64474 47640 64524 47696
rect 64460 47636 64524 47640
rect 63172 44780 63236 44844
rect 4740 44528 4804 44592
rect 4820 44528 4884 44592
rect 4900 44528 4964 44592
rect 4980 44528 5044 44592
rect 5060 44528 5124 44592
rect 5140 44528 5204 44592
rect 5220 44528 5284 44592
rect 10740 44528 10804 44592
rect 10820 44528 10884 44592
rect 10900 44528 10964 44592
rect 10980 44528 11044 44592
rect 11060 44528 11124 44592
rect 11140 44528 11204 44592
rect 11220 44528 11284 44592
rect 16740 44528 16804 44592
rect 16820 44528 16884 44592
rect 16900 44528 16964 44592
rect 16980 44528 17044 44592
rect 17060 44588 17124 44592
rect 17140 44588 17204 44592
rect 17060 44532 17100 44588
rect 17100 44532 17124 44588
rect 17140 44532 17156 44588
rect 17156 44532 17204 44588
rect 17060 44528 17124 44532
rect 17140 44528 17204 44532
rect 17220 44528 17284 44592
rect 22740 44528 22804 44592
rect 22820 44588 22884 44592
rect 22900 44588 22964 44592
rect 22820 44532 22880 44588
rect 22880 44532 22884 44588
rect 22900 44532 22936 44588
rect 22936 44532 22964 44588
rect 22820 44528 22884 44532
rect 22900 44528 22964 44532
rect 22980 44528 23044 44592
rect 23060 44528 23124 44592
rect 23140 44528 23204 44592
rect 23220 44528 23284 44592
rect 28740 44528 28804 44592
rect 28820 44528 28884 44592
rect 28900 44528 28964 44592
rect 28980 44528 29044 44592
rect 29060 44528 29124 44592
rect 29140 44528 29204 44592
rect 29220 44528 29284 44592
rect 34740 44528 34804 44592
rect 34820 44528 34884 44592
rect 34900 44528 34964 44592
rect 34980 44528 35044 44592
rect 35060 44528 35124 44592
rect 35140 44528 35204 44592
rect 35220 44528 35284 44592
rect 40740 44528 40804 44592
rect 40820 44528 40884 44592
rect 40900 44528 40964 44592
rect 40980 44528 41044 44592
rect 41060 44528 41124 44592
rect 41140 44528 41204 44592
rect 41220 44528 41284 44592
rect 46740 44528 46804 44592
rect 46820 44528 46884 44592
rect 46900 44528 46964 44592
rect 46980 44528 47044 44592
rect 47060 44528 47124 44592
rect 47140 44528 47204 44592
rect 47220 44528 47284 44592
rect 52740 44528 52804 44592
rect 52820 44528 52884 44592
rect 52900 44528 52964 44592
rect 52980 44528 53044 44592
rect 53060 44528 53124 44592
rect 53140 44528 53204 44592
rect 53220 44528 53284 44592
rect 58740 44528 58804 44592
rect 58820 44528 58884 44592
rect 58900 44528 58964 44592
rect 58980 44528 59044 44592
rect 59060 44588 59124 44592
rect 59060 44532 59104 44588
rect 59104 44532 59124 44588
rect 59060 44528 59124 44532
rect 59140 44528 59204 44592
rect 59220 44528 59284 44592
rect 64740 44528 64804 44592
rect 64820 44528 64884 44592
rect 64900 44528 64964 44592
rect 64980 44528 65044 44592
rect 65060 44528 65124 44592
rect 65140 44528 65204 44592
rect 65220 44528 65284 44592
rect 70740 44528 70804 44592
rect 70820 44528 70884 44592
rect 70900 44528 70964 44592
rect 70980 44528 71044 44592
rect 71060 44528 71124 44592
rect 71140 44528 71204 44592
rect 71220 44528 71284 44592
rect 4740 44448 4804 44512
rect 4820 44448 4884 44512
rect 4900 44448 4964 44512
rect 4980 44448 5044 44512
rect 5060 44448 5124 44512
rect 5140 44448 5204 44512
rect 5220 44448 5284 44512
rect 10740 44448 10804 44512
rect 10820 44448 10884 44512
rect 10900 44448 10964 44512
rect 10980 44448 11044 44512
rect 11060 44448 11124 44512
rect 11140 44448 11204 44512
rect 11220 44448 11284 44512
rect 16740 44448 16804 44512
rect 16820 44448 16884 44512
rect 16900 44448 16964 44512
rect 16980 44448 17044 44512
rect 17060 44508 17124 44512
rect 17140 44508 17204 44512
rect 17060 44452 17100 44508
rect 17100 44452 17124 44508
rect 17140 44452 17156 44508
rect 17156 44452 17204 44508
rect 17060 44448 17124 44452
rect 17140 44448 17204 44452
rect 17220 44448 17284 44512
rect 22740 44448 22804 44512
rect 22820 44508 22884 44512
rect 22900 44508 22964 44512
rect 22820 44452 22880 44508
rect 22880 44452 22884 44508
rect 22900 44452 22936 44508
rect 22936 44452 22964 44508
rect 22820 44448 22884 44452
rect 22900 44448 22964 44452
rect 22980 44448 23044 44512
rect 23060 44448 23124 44512
rect 23140 44448 23204 44512
rect 23220 44448 23284 44512
rect 28740 44448 28804 44512
rect 28820 44448 28884 44512
rect 28900 44448 28964 44512
rect 28980 44448 29044 44512
rect 29060 44448 29124 44512
rect 29140 44448 29204 44512
rect 29220 44448 29284 44512
rect 34740 44448 34804 44512
rect 34820 44448 34884 44512
rect 34900 44448 34964 44512
rect 34980 44448 35044 44512
rect 35060 44448 35124 44512
rect 35140 44448 35204 44512
rect 35220 44448 35284 44512
rect 40740 44448 40804 44512
rect 40820 44448 40884 44512
rect 40900 44448 40964 44512
rect 40980 44448 41044 44512
rect 41060 44448 41124 44512
rect 41140 44448 41204 44512
rect 41220 44448 41284 44512
rect 46740 44448 46804 44512
rect 46820 44448 46884 44512
rect 46900 44448 46964 44512
rect 46980 44448 47044 44512
rect 47060 44448 47124 44512
rect 47140 44448 47204 44512
rect 47220 44448 47284 44512
rect 52740 44448 52804 44512
rect 52820 44448 52884 44512
rect 52900 44448 52964 44512
rect 52980 44448 53044 44512
rect 53060 44448 53124 44512
rect 53140 44448 53204 44512
rect 53220 44448 53284 44512
rect 58740 44448 58804 44512
rect 58820 44448 58884 44512
rect 58900 44448 58964 44512
rect 58980 44448 59044 44512
rect 59060 44508 59124 44512
rect 59060 44452 59104 44508
rect 59104 44452 59124 44508
rect 59060 44448 59124 44452
rect 59140 44448 59204 44512
rect 59220 44448 59284 44512
rect 64740 44448 64804 44512
rect 64820 44448 64884 44512
rect 64900 44448 64964 44512
rect 64980 44448 65044 44512
rect 65060 44448 65124 44512
rect 65140 44448 65204 44512
rect 65220 44448 65284 44512
rect 70740 44448 70804 44512
rect 70820 44448 70884 44512
rect 70900 44448 70964 44512
rect 70980 44448 71044 44512
rect 71060 44448 71124 44512
rect 71140 44448 71204 44512
rect 71220 44448 71284 44512
rect 4740 44368 4804 44432
rect 4820 44368 4884 44432
rect 4900 44368 4964 44432
rect 4980 44368 5044 44432
rect 5060 44368 5124 44432
rect 5140 44368 5204 44432
rect 5220 44368 5284 44432
rect 10740 44368 10804 44432
rect 10820 44368 10884 44432
rect 10900 44368 10964 44432
rect 10980 44368 11044 44432
rect 11060 44368 11124 44432
rect 11140 44368 11204 44432
rect 11220 44368 11284 44432
rect 16740 44368 16804 44432
rect 16820 44368 16884 44432
rect 16900 44368 16964 44432
rect 16980 44368 17044 44432
rect 17060 44428 17124 44432
rect 17140 44428 17204 44432
rect 17060 44372 17100 44428
rect 17100 44372 17124 44428
rect 17140 44372 17156 44428
rect 17156 44372 17204 44428
rect 17060 44368 17124 44372
rect 17140 44368 17204 44372
rect 17220 44368 17284 44432
rect 22740 44368 22804 44432
rect 22820 44428 22884 44432
rect 22900 44428 22964 44432
rect 22820 44372 22880 44428
rect 22880 44372 22884 44428
rect 22900 44372 22936 44428
rect 22936 44372 22964 44428
rect 22820 44368 22884 44372
rect 22900 44368 22964 44372
rect 22980 44368 23044 44432
rect 23060 44368 23124 44432
rect 23140 44368 23204 44432
rect 23220 44368 23284 44432
rect 28740 44368 28804 44432
rect 28820 44368 28884 44432
rect 28900 44368 28964 44432
rect 28980 44368 29044 44432
rect 29060 44368 29124 44432
rect 29140 44368 29204 44432
rect 29220 44368 29284 44432
rect 34740 44368 34804 44432
rect 34820 44368 34884 44432
rect 34900 44368 34964 44432
rect 34980 44368 35044 44432
rect 35060 44368 35124 44432
rect 35140 44368 35204 44432
rect 35220 44368 35284 44432
rect 40740 44368 40804 44432
rect 40820 44368 40884 44432
rect 40900 44368 40964 44432
rect 40980 44368 41044 44432
rect 41060 44368 41124 44432
rect 41140 44368 41204 44432
rect 41220 44368 41284 44432
rect 46740 44368 46804 44432
rect 46820 44368 46884 44432
rect 46900 44368 46964 44432
rect 46980 44368 47044 44432
rect 47060 44368 47124 44432
rect 47140 44368 47204 44432
rect 47220 44368 47284 44432
rect 52740 44368 52804 44432
rect 52820 44368 52884 44432
rect 52900 44368 52964 44432
rect 52980 44368 53044 44432
rect 53060 44368 53124 44432
rect 53140 44368 53204 44432
rect 53220 44368 53284 44432
rect 58740 44368 58804 44432
rect 58820 44368 58884 44432
rect 58900 44368 58964 44432
rect 58980 44368 59044 44432
rect 59060 44428 59124 44432
rect 59060 44372 59104 44428
rect 59104 44372 59124 44428
rect 59060 44368 59124 44372
rect 59140 44368 59204 44432
rect 59220 44368 59284 44432
rect 64740 44368 64804 44432
rect 64820 44368 64884 44432
rect 64900 44368 64964 44432
rect 64980 44368 65044 44432
rect 65060 44368 65124 44432
rect 65140 44368 65204 44432
rect 65220 44368 65284 44432
rect 70740 44368 70804 44432
rect 70820 44368 70884 44432
rect 70900 44368 70964 44432
rect 70980 44368 71044 44432
rect 71060 44368 71124 44432
rect 71140 44368 71204 44432
rect 71220 44368 71284 44432
rect 4740 44288 4804 44352
rect 4820 44288 4884 44352
rect 4900 44288 4964 44352
rect 4980 44288 5044 44352
rect 5060 44288 5124 44352
rect 5140 44288 5204 44352
rect 5220 44288 5284 44352
rect 10740 44288 10804 44352
rect 10820 44288 10884 44352
rect 10900 44288 10964 44352
rect 10980 44288 11044 44352
rect 11060 44288 11124 44352
rect 11140 44288 11204 44352
rect 11220 44288 11284 44352
rect 16740 44288 16804 44352
rect 16820 44288 16884 44352
rect 16900 44288 16964 44352
rect 16980 44288 17044 44352
rect 17060 44348 17124 44352
rect 17140 44348 17204 44352
rect 17060 44292 17100 44348
rect 17100 44292 17124 44348
rect 17140 44292 17156 44348
rect 17156 44292 17204 44348
rect 17060 44288 17124 44292
rect 17140 44288 17204 44292
rect 17220 44288 17284 44352
rect 22740 44288 22804 44352
rect 22820 44348 22884 44352
rect 22900 44348 22964 44352
rect 22820 44292 22880 44348
rect 22880 44292 22884 44348
rect 22900 44292 22936 44348
rect 22936 44292 22964 44348
rect 22820 44288 22884 44292
rect 22900 44288 22964 44292
rect 22980 44288 23044 44352
rect 23060 44288 23124 44352
rect 23140 44288 23204 44352
rect 23220 44288 23284 44352
rect 28740 44288 28804 44352
rect 28820 44288 28884 44352
rect 28900 44288 28964 44352
rect 28980 44288 29044 44352
rect 29060 44288 29124 44352
rect 29140 44288 29204 44352
rect 29220 44288 29284 44352
rect 34740 44288 34804 44352
rect 34820 44288 34884 44352
rect 34900 44288 34964 44352
rect 34980 44288 35044 44352
rect 35060 44288 35124 44352
rect 35140 44288 35204 44352
rect 35220 44288 35284 44352
rect 40740 44288 40804 44352
rect 40820 44288 40884 44352
rect 40900 44288 40964 44352
rect 40980 44288 41044 44352
rect 41060 44288 41124 44352
rect 41140 44288 41204 44352
rect 41220 44288 41284 44352
rect 46740 44288 46804 44352
rect 46820 44288 46884 44352
rect 46900 44288 46964 44352
rect 46980 44288 47044 44352
rect 47060 44288 47124 44352
rect 47140 44288 47204 44352
rect 47220 44288 47284 44352
rect 52740 44288 52804 44352
rect 52820 44288 52884 44352
rect 52900 44288 52964 44352
rect 52980 44288 53044 44352
rect 53060 44288 53124 44352
rect 53140 44288 53204 44352
rect 53220 44288 53284 44352
rect 58740 44288 58804 44352
rect 58820 44288 58884 44352
rect 58900 44288 58964 44352
rect 58980 44288 59044 44352
rect 59060 44348 59124 44352
rect 59060 44292 59104 44348
rect 59104 44292 59124 44348
rect 59060 44288 59124 44292
rect 59140 44288 59204 44352
rect 59220 44288 59284 44352
rect 64740 44288 64804 44352
rect 64820 44288 64884 44352
rect 64900 44288 64964 44352
rect 64980 44288 65044 44352
rect 65060 44288 65124 44352
rect 65140 44288 65204 44352
rect 65220 44288 65284 44352
rect 70740 44288 70804 44352
rect 70820 44288 70884 44352
rect 70900 44288 70964 44352
rect 70980 44288 71044 44352
rect 71060 44288 71124 44352
rect 71140 44288 71204 44352
rect 71220 44288 71284 44352
rect 63908 43284 63972 43348
rect 1740 42176 1804 42240
rect 1820 42176 1884 42240
rect 1900 42176 1964 42240
rect 1980 42176 2044 42240
rect 2060 42176 2124 42240
rect 2140 42236 2204 42240
rect 2220 42236 2284 42240
rect 2140 42180 2184 42236
rect 2184 42180 2204 42236
rect 2220 42180 2240 42236
rect 2240 42180 2264 42236
rect 2264 42180 2284 42236
rect 2140 42176 2204 42180
rect 2220 42176 2284 42180
rect 7740 42176 7804 42240
rect 7820 42176 7884 42240
rect 7900 42176 7964 42240
rect 7980 42176 8044 42240
rect 8060 42176 8124 42240
rect 8140 42176 8204 42240
rect 8220 42236 8284 42240
rect 8220 42180 8283 42236
rect 8283 42180 8284 42236
rect 8220 42176 8284 42180
rect 13740 42176 13804 42240
rect 13820 42176 13884 42240
rect 13900 42176 13964 42240
rect 13980 42176 14044 42240
rect 14060 42236 14124 42240
rect 14060 42180 14063 42236
rect 14063 42180 14119 42236
rect 14119 42180 14124 42236
rect 14060 42176 14124 42180
rect 14140 42176 14204 42240
rect 14220 42176 14284 42240
rect 19740 42176 19804 42240
rect 19820 42236 19884 42240
rect 19820 42180 19843 42236
rect 19843 42180 19884 42236
rect 19820 42176 19884 42180
rect 19900 42176 19964 42240
rect 19980 42176 20044 42240
rect 20060 42176 20124 42240
rect 20140 42176 20204 42240
rect 20220 42176 20284 42240
rect 25740 42176 25804 42240
rect 25820 42176 25884 42240
rect 25900 42176 25964 42240
rect 25980 42176 26044 42240
rect 26060 42176 26124 42240
rect 26140 42176 26204 42240
rect 26220 42176 26284 42240
rect 31740 42176 31804 42240
rect 31820 42176 31884 42240
rect 31900 42176 31964 42240
rect 31980 42176 32044 42240
rect 32060 42176 32124 42240
rect 32140 42176 32204 42240
rect 32220 42176 32284 42240
rect 37740 42176 37804 42240
rect 37820 42176 37884 42240
rect 37900 42176 37964 42240
rect 37980 42176 38044 42240
rect 38060 42176 38124 42240
rect 38140 42176 38204 42240
rect 38220 42176 38284 42240
rect 43740 42176 43804 42240
rect 43820 42176 43884 42240
rect 43900 42176 43964 42240
rect 43980 42176 44044 42240
rect 44060 42176 44124 42240
rect 44140 42176 44204 42240
rect 44220 42176 44284 42240
rect 49740 42236 49804 42240
rect 49740 42180 49742 42236
rect 49742 42180 49798 42236
rect 49798 42180 49804 42236
rect 49740 42176 49804 42180
rect 49820 42176 49884 42240
rect 49900 42176 49964 42240
rect 49980 42176 50044 42240
rect 50060 42176 50124 42240
rect 50140 42176 50204 42240
rect 50220 42176 50284 42240
rect 55740 42176 55804 42240
rect 55820 42176 55884 42240
rect 55900 42176 55964 42240
rect 55980 42176 56044 42240
rect 56060 42176 56124 42240
rect 56140 42176 56204 42240
rect 56220 42176 56284 42240
rect 61740 42176 61804 42240
rect 61820 42176 61884 42240
rect 61900 42176 61964 42240
rect 61980 42176 62044 42240
rect 62060 42176 62124 42240
rect 62140 42176 62204 42240
rect 62220 42176 62284 42240
rect 67740 42176 67804 42240
rect 67820 42176 67884 42240
rect 67900 42176 67964 42240
rect 67980 42176 68044 42240
rect 68060 42176 68124 42240
rect 68140 42176 68204 42240
rect 68220 42176 68284 42240
rect 73740 42176 73804 42240
rect 73820 42176 73884 42240
rect 73900 42176 73964 42240
rect 73980 42176 74044 42240
rect 74060 42176 74124 42240
rect 74140 42176 74204 42240
rect 74220 42176 74284 42240
rect 1740 42096 1804 42160
rect 1820 42096 1884 42160
rect 1900 42096 1964 42160
rect 1980 42096 2044 42160
rect 2060 42096 2124 42160
rect 2140 42156 2204 42160
rect 2220 42156 2284 42160
rect 2140 42100 2184 42156
rect 2184 42100 2204 42156
rect 2220 42100 2240 42156
rect 2240 42100 2264 42156
rect 2264 42100 2284 42156
rect 2140 42096 2204 42100
rect 2220 42096 2284 42100
rect 7740 42096 7804 42160
rect 7820 42096 7884 42160
rect 7900 42096 7964 42160
rect 7980 42096 8044 42160
rect 8060 42096 8124 42160
rect 8140 42096 8204 42160
rect 8220 42156 8284 42160
rect 8220 42100 8283 42156
rect 8283 42100 8284 42156
rect 8220 42096 8284 42100
rect 13740 42096 13804 42160
rect 13820 42096 13884 42160
rect 13900 42096 13964 42160
rect 13980 42096 14044 42160
rect 14060 42156 14124 42160
rect 14060 42100 14063 42156
rect 14063 42100 14119 42156
rect 14119 42100 14124 42156
rect 14060 42096 14124 42100
rect 14140 42096 14204 42160
rect 14220 42096 14284 42160
rect 19740 42096 19804 42160
rect 19820 42156 19884 42160
rect 19820 42100 19843 42156
rect 19843 42100 19884 42156
rect 19820 42096 19884 42100
rect 19900 42096 19964 42160
rect 19980 42096 20044 42160
rect 20060 42096 20124 42160
rect 20140 42096 20204 42160
rect 20220 42096 20284 42160
rect 25740 42096 25804 42160
rect 25820 42096 25884 42160
rect 25900 42096 25964 42160
rect 25980 42096 26044 42160
rect 26060 42096 26124 42160
rect 26140 42096 26204 42160
rect 26220 42096 26284 42160
rect 31740 42096 31804 42160
rect 31820 42096 31884 42160
rect 31900 42096 31964 42160
rect 31980 42096 32044 42160
rect 32060 42096 32124 42160
rect 32140 42096 32204 42160
rect 32220 42096 32284 42160
rect 37740 42096 37804 42160
rect 37820 42096 37884 42160
rect 37900 42096 37964 42160
rect 37980 42096 38044 42160
rect 38060 42096 38124 42160
rect 38140 42096 38204 42160
rect 38220 42096 38284 42160
rect 43740 42096 43804 42160
rect 43820 42096 43884 42160
rect 43900 42096 43964 42160
rect 43980 42096 44044 42160
rect 44060 42096 44124 42160
rect 44140 42096 44204 42160
rect 44220 42096 44284 42160
rect 49740 42156 49804 42160
rect 49740 42100 49742 42156
rect 49742 42100 49798 42156
rect 49798 42100 49804 42156
rect 49740 42096 49804 42100
rect 49820 42096 49884 42160
rect 49900 42096 49964 42160
rect 49980 42096 50044 42160
rect 50060 42096 50124 42160
rect 50140 42096 50204 42160
rect 50220 42096 50284 42160
rect 55740 42096 55804 42160
rect 55820 42096 55884 42160
rect 55900 42096 55964 42160
rect 55980 42096 56044 42160
rect 56060 42096 56124 42160
rect 56140 42096 56204 42160
rect 56220 42096 56284 42160
rect 61740 42096 61804 42160
rect 61820 42096 61884 42160
rect 61900 42096 61964 42160
rect 61980 42096 62044 42160
rect 62060 42096 62124 42160
rect 62140 42096 62204 42160
rect 62220 42096 62284 42160
rect 67740 42096 67804 42160
rect 67820 42096 67884 42160
rect 67900 42096 67964 42160
rect 67980 42096 68044 42160
rect 68060 42096 68124 42160
rect 68140 42096 68204 42160
rect 68220 42096 68284 42160
rect 73740 42096 73804 42160
rect 73820 42096 73884 42160
rect 73900 42096 73964 42160
rect 73980 42096 74044 42160
rect 74060 42096 74124 42160
rect 74140 42096 74204 42160
rect 74220 42096 74284 42160
rect 1740 42016 1804 42080
rect 1820 42016 1884 42080
rect 1900 42016 1964 42080
rect 1980 42016 2044 42080
rect 2060 42016 2124 42080
rect 2140 42076 2204 42080
rect 2220 42076 2284 42080
rect 2140 42020 2184 42076
rect 2184 42020 2204 42076
rect 2220 42020 2240 42076
rect 2240 42020 2264 42076
rect 2264 42020 2284 42076
rect 2140 42016 2204 42020
rect 2220 42016 2284 42020
rect 7740 42016 7804 42080
rect 7820 42016 7884 42080
rect 7900 42016 7964 42080
rect 7980 42016 8044 42080
rect 8060 42016 8124 42080
rect 8140 42016 8204 42080
rect 8220 42076 8284 42080
rect 8220 42020 8283 42076
rect 8283 42020 8284 42076
rect 8220 42016 8284 42020
rect 13740 42016 13804 42080
rect 13820 42016 13884 42080
rect 13900 42016 13964 42080
rect 13980 42016 14044 42080
rect 14060 42076 14124 42080
rect 14060 42020 14063 42076
rect 14063 42020 14119 42076
rect 14119 42020 14124 42076
rect 14060 42016 14124 42020
rect 14140 42016 14204 42080
rect 14220 42016 14284 42080
rect 19740 42016 19804 42080
rect 19820 42076 19884 42080
rect 19820 42020 19843 42076
rect 19843 42020 19884 42076
rect 19820 42016 19884 42020
rect 19900 42016 19964 42080
rect 19980 42016 20044 42080
rect 20060 42016 20124 42080
rect 20140 42016 20204 42080
rect 20220 42016 20284 42080
rect 25740 42016 25804 42080
rect 25820 42016 25884 42080
rect 25900 42016 25964 42080
rect 25980 42016 26044 42080
rect 26060 42016 26124 42080
rect 26140 42016 26204 42080
rect 26220 42016 26284 42080
rect 31740 42016 31804 42080
rect 31820 42016 31884 42080
rect 31900 42016 31964 42080
rect 31980 42016 32044 42080
rect 32060 42016 32124 42080
rect 32140 42016 32204 42080
rect 32220 42016 32284 42080
rect 37740 42016 37804 42080
rect 37820 42016 37884 42080
rect 37900 42016 37964 42080
rect 37980 42016 38044 42080
rect 38060 42016 38124 42080
rect 38140 42016 38204 42080
rect 38220 42016 38284 42080
rect 43740 42016 43804 42080
rect 43820 42016 43884 42080
rect 43900 42016 43964 42080
rect 43980 42016 44044 42080
rect 44060 42016 44124 42080
rect 44140 42016 44204 42080
rect 44220 42016 44284 42080
rect 49740 42076 49804 42080
rect 49740 42020 49742 42076
rect 49742 42020 49798 42076
rect 49798 42020 49804 42076
rect 49740 42016 49804 42020
rect 49820 42016 49884 42080
rect 49900 42016 49964 42080
rect 49980 42016 50044 42080
rect 50060 42016 50124 42080
rect 50140 42016 50204 42080
rect 50220 42016 50284 42080
rect 55740 42016 55804 42080
rect 55820 42016 55884 42080
rect 55900 42016 55964 42080
rect 55980 42016 56044 42080
rect 56060 42016 56124 42080
rect 56140 42016 56204 42080
rect 56220 42016 56284 42080
rect 61740 42016 61804 42080
rect 61820 42016 61884 42080
rect 61900 42016 61964 42080
rect 61980 42016 62044 42080
rect 62060 42016 62124 42080
rect 62140 42016 62204 42080
rect 62220 42016 62284 42080
rect 67740 42016 67804 42080
rect 67820 42016 67884 42080
rect 67900 42016 67964 42080
rect 67980 42016 68044 42080
rect 68060 42016 68124 42080
rect 68140 42016 68204 42080
rect 68220 42016 68284 42080
rect 73740 42016 73804 42080
rect 73820 42016 73884 42080
rect 73900 42016 73964 42080
rect 73980 42016 74044 42080
rect 74060 42016 74124 42080
rect 74140 42016 74204 42080
rect 74220 42016 74284 42080
rect 1740 41936 1804 42000
rect 1820 41936 1884 42000
rect 1900 41936 1964 42000
rect 1980 41936 2044 42000
rect 2060 41936 2124 42000
rect 2140 41996 2204 42000
rect 2220 41996 2284 42000
rect 2140 41940 2184 41996
rect 2184 41940 2204 41996
rect 2220 41940 2240 41996
rect 2240 41940 2264 41996
rect 2264 41940 2284 41996
rect 2140 41936 2204 41940
rect 2220 41936 2284 41940
rect 7740 41936 7804 42000
rect 7820 41936 7884 42000
rect 7900 41936 7964 42000
rect 7980 41936 8044 42000
rect 8060 41936 8124 42000
rect 8140 41936 8204 42000
rect 8220 41996 8284 42000
rect 8220 41940 8283 41996
rect 8283 41940 8284 41996
rect 8220 41936 8284 41940
rect 13740 41936 13804 42000
rect 13820 41936 13884 42000
rect 13900 41936 13964 42000
rect 13980 41936 14044 42000
rect 14060 41996 14124 42000
rect 14060 41940 14063 41996
rect 14063 41940 14119 41996
rect 14119 41940 14124 41996
rect 14060 41936 14124 41940
rect 14140 41936 14204 42000
rect 14220 41936 14284 42000
rect 19740 41936 19804 42000
rect 19820 41996 19884 42000
rect 19820 41940 19843 41996
rect 19843 41940 19884 41996
rect 19820 41936 19884 41940
rect 19900 41936 19964 42000
rect 19980 41936 20044 42000
rect 20060 41936 20124 42000
rect 20140 41936 20204 42000
rect 20220 41936 20284 42000
rect 25740 41936 25804 42000
rect 25820 41936 25884 42000
rect 25900 41936 25964 42000
rect 25980 41936 26044 42000
rect 26060 41936 26124 42000
rect 26140 41936 26204 42000
rect 26220 41936 26284 42000
rect 31740 41936 31804 42000
rect 31820 41936 31884 42000
rect 31900 41936 31964 42000
rect 31980 41936 32044 42000
rect 32060 41936 32124 42000
rect 32140 41936 32204 42000
rect 32220 41936 32284 42000
rect 37740 41936 37804 42000
rect 37820 41936 37884 42000
rect 37900 41936 37964 42000
rect 37980 41936 38044 42000
rect 38060 41936 38124 42000
rect 38140 41936 38204 42000
rect 38220 41936 38284 42000
rect 43740 41936 43804 42000
rect 43820 41936 43884 42000
rect 43900 41936 43964 42000
rect 43980 41936 44044 42000
rect 44060 41936 44124 42000
rect 44140 41936 44204 42000
rect 44220 41936 44284 42000
rect 49740 41996 49804 42000
rect 49740 41940 49742 41996
rect 49742 41940 49798 41996
rect 49798 41940 49804 41996
rect 49740 41936 49804 41940
rect 49820 41936 49884 42000
rect 49900 41936 49964 42000
rect 49980 41936 50044 42000
rect 50060 41936 50124 42000
rect 50140 41936 50204 42000
rect 50220 41936 50284 42000
rect 55740 41936 55804 42000
rect 55820 41936 55884 42000
rect 55900 41936 55964 42000
rect 55980 41936 56044 42000
rect 56060 41936 56124 42000
rect 56140 41936 56204 42000
rect 56220 41936 56284 42000
rect 61740 41936 61804 42000
rect 61820 41936 61884 42000
rect 61900 41936 61964 42000
rect 61980 41936 62044 42000
rect 62060 41936 62124 42000
rect 62140 41936 62204 42000
rect 62220 41936 62284 42000
rect 67740 41936 67804 42000
rect 67820 41936 67884 42000
rect 67900 41936 67964 42000
rect 67980 41936 68044 42000
rect 68060 41936 68124 42000
rect 68140 41936 68204 42000
rect 68220 41936 68284 42000
rect 73740 41936 73804 42000
rect 73820 41936 73884 42000
rect 73900 41936 73964 42000
rect 73980 41936 74044 42000
rect 74060 41936 74124 42000
rect 74140 41936 74204 42000
rect 74220 41936 74284 42000
rect 65748 40836 65812 40900
rect 65932 38660 65996 38724
rect 4740 34528 4804 34592
rect 4820 34528 4884 34592
rect 4900 34528 4964 34592
rect 4980 34528 5044 34592
rect 5060 34528 5124 34592
rect 5140 34528 5204 34592
rect 5220 34528 5284 34592
rect 10740 34528 10804 34592
rect 10820 34528 10884 34592
rect 10900 34528 10964 34592
rect 10980 34528 11044 34592
rect 11060 34528 11124 34592
rect 11140 34528 11204 34592
rect 11220 34528 11284 34592
rect 16740 34528 16804 34592
rect 16820 34528 16884 34592
rect 16900 34528 16964 34592
rect 16980 34528 17044 34592
rect 17060 34588 17124 34592
rect 17140 34588 17204 34592
rect 17060 34532 17100 34588
rect 17100 34532 17124 34588
rect 17140 34532 17156 34588
rect 17156 34532 17204 34588
rect 17060 34528 17124 34532
rect 17140 34528 17204 34532
rect 17220 34528 17284 34592
rect 22740 34528 22804 34592
rect 22820 34588 22884 34592
rect 22900 34588 22964 34592
rect 22820 34532 22880 34588
rect 22880 34532 22884 34588
rect 22900 34532 22936 34588
rect 22936 34532 22964 34588
rect 22820 34528 22884 34532
rect 22900 34528 22964 34532
rect 22980 34528 23044 34592
rect 23060 34528 23124 34592
rect 23140 34528 23204 34592
rect 23220 34528 23284 34592
rect 28740 34528 28804 34592
rect 28820 34528 28884 34592
rect 28900 34528 28964 34592
rect 28980 34528 29044 34592
rect 29060 34528 29124 34592
rect 29140 34528 29204 34592
rect 29220 34528 29284 34592
rect 34740 34528 34804 34592
rect 34820 34528 34884 34592
rect 34900 34528 34964 34592
rect 34980 34528 35044 34592
rect 35060 34528 35124 34592
rect 35140 34528 35204 34592
rect 35220 34528 35284 34592
rect 40740 34528 40804 34592
rect 40820 34528 40884 34592
rect 40900 34528 40964 34592
rect 40980 34528 41044 34592
rect 41060 34528 41124 34592
rect 41140 34528 41204 34592
rect 41220 34528 41284 34592
rect 46740 34528 46804 34592
rect 46820 34528 46884 34592
rect 46900 34528 46964 34592
rect 46980 34528 47044 34592
rect 47060 34528 47124 34592
rect 47140 34528 47204 34592
rect 47220 34528 47284 34592
rect 52740 34528 52804 34592
rect 52820 34528 52884 34592
rect 52900 34528 52964 34592
rect 52980 34528 53044 34592
rect 53060 34528 53124 34592
rect 53140 34528 53204 34592
rect 53220 34528 53284 34592
rect 58740 34528 58804 34592
rect 58820 34528 58884 34592
rect 58900 34528 58964 34592
rect 58980 34528 59044 34592
rect 59060 34588 59124 34592
rect 59060 34532 59104 34588
rect 59104 34532 59124 34588
rect 59060 34528 59124 34532
rect 59140 34528 59204 34592
rect 59220 34528 59284 34592
rect 64740 34528 64804 34592
rect 64820 34528 64884 34592
rect 64900 34528 64964 34592
rect 64980 34528 65044 34592
rect 65060 34528 65124 34592
rect 65140 34528 65204 34592
rect 65220 34528 65284 34592
rect 70740 34528 70804 34592
rect 70820 34528 70884 34592
rect 70900 34528 70964 34592
rect 70980 34528 71044 34592
rect 71060 34528 71124 34592
rect 71140 34528 71204 34592
rect 71220 34528 71284 34592
rect 4740 34448 4804 34512
rect 4820 34448 4884 34512
rect 4900 34448 4964 34512
rect 4980 34448 5044 34512
rect 5060 34448 5124 34512
rect 5140 34448 5204 34512
rect 5220 34448 5284 34512
rect 10740 34448 10804 34512
rect 10820 34448 10884 34512
rect 10900 34448 10964 34512
rect 10980 34448 11044 34512
rect 11060 34448 11124 34512
rect 11140 34448 11204 34512
rect 11220 34448 11284 34512
rect 16740 34448 16804 34512
rect 16820 34448 16884 34512
rect 16900 34448 16964 34512
rect 16980 34448 17044 34512
rect 17060 34508 17124 34512
rect 17140 34508 17204 34512
rect 17060 34452 17100 34508
rect 17100 34452 17124 34508
rect 17140 34452 17156 34508
rect 17156 34452 17204 34508
rect 17060 34448 17124 34452
rect 17140 34448 17204 34452
rect 17220 34448 17284 34512
rect 22740 34448 22804 34512
rect 22820 34508 22884 34512
rect 22900 34508 22964 34512
rect 22820 34452 22880 34508
rect 22880 34452 22884 34508
rect 22900 34452 22936 34508
rect 22936 34452 22964 34508
rect 22820 34448 22884 34452
rect 22900 34448 22964 34452
rect 22980 34448 23044 34512
rect 23060 34448 23124 34512
rect 23140 34448 23204 34512
rect 23220 34448 23284 34512
rect 28740 34448 28804 34512
rect 28820 34448 28884 34512
rect 28900 34448 28964 34512
rect 28980 34448 29044 34512
rect 29060 34448 29124 34512
rect 29140 34448 29204 34512
rect 29220 34448 29284 34512
rect 34740 34448 34804 34512
rect 34820 34448 34884 34512
rect 34900 34448 34964 34512
rect 34980 34448 35044 34512
rect 35060 34448 35124 34512
rect 35140 34448 35204 34512
rect 35220 34448 35284 34512
rect 40740 34448 40804 34512
rect 40820 34448 40884 34512
rect 40900 34448 40964 34512
rect 40980 34448 41044 34512
rect 41060 34448 41124 34512
rect 41140 34448 41204 34512
rect 41220 34448 41284 34512
rect 46740 34448 46804 34512
rect 46820 34448 46884 34512
rect 46900 34448 46964 34512
rect 46980 34448 47044 34512
rect 47060 34448 47124 34512
rect 47140 34448 47204 34512
rect 47220 34448 47284 34512
rect 52740 34448 52804 34512
rect 52820 34448 52884 34512
rect 52900 34448 52964 34512
rect 52980 34448 53044 34512
rect 53060 34448 53124 34512
rect 53140 34448 53204 34512
rect 53220 34448 53284 34512
rect 58740 34448 58804 34512
rect 58820 34448 58884 34512
rect 58900 34448 58964 34512
rect 58980 34448 59044 34512
rect 59060 34508 59124 34512
rect 59060 34452 59104 34508
rect 59104 34452 59124 34508
rect 59060 34448 59124 34452
rect 59140 34448 59204 34512
rect 59220 34448 59284 34512
rect 64740 34448 64804 34512
rect 64820 34448 64884 34512
rect 64900 34448 64964 34512
rect 64980 34448 65044 34512
rect 65060 34448 65124 34512
rect 65140 34448 65204 34512
rect 65220 34448 65284 34512
rect 70740 34448 70804 34512
rect 70820 34448 70884 34512
rect 70900 34448 70964 34512
rect 70980 34448 71044 34512
rect 71060 34448 71124 34512
rect 71140 34448 71204 34512
rect 71220 34448 71284 34512
rect 4740 34368 4804 34432
rect 4820 34368 4884 34432
rect 4900 34368 4964 34432
rect 4980 34368 5044 34432
rect 5060 34368 5124 34432
rect 5140 34368 5204 34432
rect 5220 34368 5284 34432
rect 10740 34368 10804 34432
rect 10820 34368 10884 34432
rect 10900 34368 10964 34432
rect 10980 34368 11044 34432
rect 11060 34368 11124 34432
rect 11140 34368 11204 34432
rect 11220 34368 11284 34432
rect 16740 34368 16804 34432
rect 16820 34368 16884 34432
rect 16900 34368 16964 34432
rect 16980 34368 17044 34432
rect 17060 34428 17124 34432
rect 17140 34428 17204 34432
rect 17060 34372 17100 34428
rect 17100 34372 17124 34428
rect 17140 34372 17156 34428
rect 17156 34372 17204 34428
rect 17060 34368 17124 34372
rect 17140 34368 17204 34372
rect 17220 34368 17284 34432
rect 22740 34368 22804 34432
rect 22820 34428 22884 34432
rect 22900 34428 22964 34432
rect 22820 34372 22880 34428
rect 22880 34372 22884 34428
rect 22900 34372 22936 34428
rect 22936 34372 22964 34428
rect 22820 34368 22884 34372
rect 22900 34368 22964 34372
rect 22980 34368 23044 34432
rect 23060 34368 23124 34432
rect 23140 34368 23204 34432
rect 23220 34368 23284 34432
rect 28740 34368 28804 34432
rect 28820 34368 28884 34432
rect 28900 34368 28964 34432
rect 28980 34368 29044 34432
rect 29060 34368 29124 34432
rect 29140 34368 29204 34432
rect 29220 34368 29284 34432
rect 34740 34368 34804 34432
rect 34820 34368 34884 34432
rect 34900 34368 34964 34432
rect 34980 34368 35044 34432
rect 35060 34368 35124 34432
rect 35140 34368 35204 34432
rect 35220 34368 35284 34432
rect 40740 34368 40804 34432
rect 40820 34368 40884 34432
rect 40900 34368 40964 34432
rect 40980 34368 41044 34432
rect 41060 34368 41124 34432
rect 41140 34368 41204 34432
rect 41220 34368 41284 34432
rect 46740 34368 46804 34432
rect 46820 34368 46884 34432
rect 46900 34368 46964 34432
rect 46980 34368 47044 34432
rect 47060 34368 47124 34432
rect 47140 34368 47204 34432
rect 47220 34368 47284 34432
rect 52740 34368 52804 34432
rect 52820 34368 52884 34432
rect 52900 34368 52964 34432
rect 52980 34368 53044 34432
rect 53060 34368 53124 34432
rect 53140 34368 53204 34432
rect 53220 34368 53284 34432
rect 58740 34368 58804 34432
rect 58820 34368 58884 34432
rect 58900 34368 58964 34432
rect 58980 34368 59044 34432
rect 59060 34428 59124 34432
rect 59060 34372 59104 34428
rect 59104 34372 59124 34428
rect 59060 34368 59124 34372
rect 59140 34368 59204 34432
rect 59220 34368 59284 34432
rect 64740 34368 64804 34432
rect 64820 34368 64884 34432
rect 64900 34368 64964 34432
rect 64980 34368 65044 34432
rect 65060 34368 65124 34432
rect 65140 34368 65204 34432
rect 65220 34368 65284 34432
rect 70740 34368 70804 34432
rect 70820 34368 70884 34432
rect 70900 34368 70964 34432
rect 70980 34368 71044 34432
rect 71060 34368 71124 34432
rect 71140 34368 71204 34432
rect 71220 34368 71284 34432
rect 4740 34288 4804 34352
rect 4820 34288 4884 34352
rect 4900 34288 4964 34352
rect 4980 34288 5044 34352
rect 5060 34288 5124 34352
rect 5140 34288 5204 34352
rect 5220 34288 5284 34352
rect 10740 34288 10804 34352
rect 10820 34288 10884 34352
rect 10900 34288 10964 34352
rect 10980 34288 11044 34352
rect 11060 34288 11124 34352
rect 11140 34288 11204 34352
rect 11220 34288 11284 34352
rect 16740 34288 16804 34352
rect 16820 34288 16884 34352
rect 16900 34288 16964 34352
rect 16980 34288 17044 34352
rect 17060 34348 17124 34352
rect 17140 34348 17204 34352
rect 17060 34292 17100 34348
rect 17100 34292 17124 34348
rect 17140 34292 17156 34348
rect 17156 34292 17204 34348
rect 17060 34288 17124 34292
rect 17140 34288 17204 34292
rect 17220 34288 17284 34352
rect 22740 34288 22804 34352
rect 22820 34348 22884 34352
rect 22900 34348 22964 34352
rect 22820 34292 22880 34348
rect 22880 34292 22884 34348
rect 22900 34292 22936 34348
rect 22936 34292 22964 34348
rect 22820 34288 22884 34292
rect 22900 34288 22964 34292
rect 22980 34288 23044 34352
rect 23060 34288 23124 34352
rect 23140 34288 23204 34352
rect 23220 34288 23284 34352
rect 28740 34288 28804 34352
rect 28820 34288 28884 34352
rect 28900 34288 28964 34352
rect 28980 34288 29044 34352
rect 29060 34288 29124 34352
rect 29140 34288 29204 34352
rect 29220 34288 29284 34352
rect 34740 34288 34804 34352
rect 34820 34288 34884 34352
rect 34900 34288 34964 34352
rect 34980 34288 35044 34352
rect 35060 34288 35124 34352
rect 35140 34288 35204 34352
rect 35220 34288 35284 34352
rect 40740 34288 40804 34352
rect 40820 34288 40884 34352
rect 40900 34288 40964 34352
rect 40980 34288 41044 34352
rect 41060 34288 41124 34352
rect 41140 34288 41204 34352
rect 41220 34288 41284 34352
rect 46740 34288 46804 34352
rect 46820 34288 46884 34352
rect 46900 34288 46964 34352
rect 46980 34288 47044 34352
rect 47060 34288 47124 34352
rect 47140 34288 47204 34352
rect 47220 34288 47284 34352
rect 52740 34288 52804 34352
rect 52820 34288 52884 34352
rect 52900 34288 52964 34352
rect 52980 34288 53044 34352
rect 53060 34288 53124 34352
rect 53140 34288 53204 34352
rect 53220 34288 53284 34352
rect 58740 34288 58804 34352
rect 58820 34288 58884 34352
rect 58900 34288 58964 34352
rect 58980 34288 59044 34352
rect 59060 34348 59124 34352
rect 59060 34292 59104 34348
rect 59104 34292 59124 34348
rect 59060 34288 59124 34292
rect 59140 34288 59204 34352
rect 59220 34288 59284 34352
rect 64740 34288 64804 34352
rect 64820 34288 64884 34352
rect 64900 34288 64964 34352
rect 64980 34288 65044 34352
rect 65060 34288 65124 34352
rect 65140 34288 65204 34352
rect 65220 34288 65284 34352
rect 70740 34288 70804 34352
rect 70820 34288 70884 34352
rect 70900 34288 70964 34352
rect 70980 34288 71044 34352
rect 71060 34288 71124 34352
rect 71140 34288 71204 34352
rect 71220 34288 71284 34352
rect 68508 33220 68572 33284
rect 1740 32176 1804 32240
rect 1820 32176 1884 32240
rect 1900 32176 1964 32240
rect 1980 32176 2044 32240
rect 2060 32176 2124 32240
rect 2140 32236 2204 32240
rect 2220 32236 2284 32240
rect 2140 32180 2184 32236
rect 2184 32180 2204 32236
rect 2220 32180 2240 32236
rect 2240 32180 2264 32236
rect 2264 32180 2284 32236
rect 2140 32176 2204 32180
rect 2220 32176 2284 32180
rect 7740 32176 7804 32240
rect 7820 32176 7884 32240
rect 7900 32176 7964 32240
rect 7980 32176 8044 32240
rect 8060 32176 8124 32240
rect 8140 32176 8204 32240
rect 8220 32236 8284 32240
rect 8220 32180 8283 32236
rect 8283 32180 8284 32236
rect 8220 32176 8284 32180
rect 13740 32176 13804 32240
rect 13820 32176 13884 32240
rect 13900 32176 13964 32240
rect 13980 32176 14044 32240
rect 14060 32236 14124 32240
rect 14060 32180 14063 32236
rect 14063 32180 14119 32236
rect 14119 32180 14124 32236
rect 14060 32176 14124 32180
rect 14140 32176 14204 32240
rect 14220 32176 14284 32240
rect 19740 32176 19804 32240
rect 19820 32236 19884 32240
rect 19820 32180 19843 32236
rect 19843 32180 19884 32236
rect 19820 32176 19884 32180
rect 19900 32176 19964 32240
rect 19980 32176 20044 32240
rect 20060 32176 20124 32240
rect 20140 32176 20204 32240
rect 20220 32176 20284 32240
rect 25740 32176 25804 32240
rect 25820 32176 25884 32240
rect 25900 32176 25964 32240
rect 25980 32176 26044 32240
rect 26060 32176 26124 32240
rect 26140 32176 26204 32240
rect 26220 32176 26284 32240
rect 31740 32176 31804 32240
rect 31820 32176 31884 32240
rect 31900 32176 31964 32240
rect 31980 32176 32044 32240
rect 32060 32176 32124 32240
rect 32140 32176 32204 32240
rect 32220 32176 32284 32240
rect 37740 32176 37804 32240
rect 37820 32176 37884 32240
rect 37900 32176 37964 32240
rect 37980 32176 38044 32240
rect 38060 32176 38124 32240
rect 38140 32176 38204 32240
rect 38220 32176 38284 32240
rect 43740 32176 43804 32240
rect 43820 32176 43884 32240
rect 43900 32176 43964 32240
rect 43980 32176 44044 32240
rect 44060 32176 44124 32240
rect 44140 32176 44204 32240
rect 44220 32176 44284 32240
rect 49740 32236 49804 32240
rect 49740 32180 49742 32236
rect 49742 32180 49798 32236
rect 49798 32180 49804 32236
rect 49740 32176 49804 32180
rect 49820 32176 49884 32240
rect 49900 32176 49964 32240
rect 49980 32176 50044 32240
rect 50060 32176 50124 32240
rect 50140 32176 50204 32240
rect 50220 32176 50284 32240
rect 55740 32176 55804 32240
rect 55820 32176 55884 32240
rect 55900 32176 55964 32240
rect 55980 32176 56044 32240
rect 56060 32176 56124 32240
rect 56140 32176 56204 32240
rect 56220 32176 56284 32240
rect 61740 32176 61804 32240
rect 61820 32176 61884 32240
rect 61900 32176 61964 32240
rect 61980 32176 62044 32240
rect 62060 32176 62124 32240
rect 62140 32176 62204 32240
rect 62220 32176 62284 32240
rect 67740 32176 67804 32240
rect 67820 32176 67884 32240
rect 67900 32176 67964 32240
rect 67980 32176 68044 32240
rect 68060 32176 68124 32240
rect 68140 32176 68204 32240
rect 68220 32176 68284 32240
rect 73740 32176 73804 32240
rect 73820 32176 73884 32240
rect 73900 32176 73964 32240
rect 73980 32176 74044 32240
rect 74060 32176 74124 32240
rect 74140 32176 74204 32240
rect 74220 32176 74284 32240
rect 1740 32096 1804 32160
rect 1820 32096 1884 32160
rect 1900 32096 1964 32160
rect 1980 32096 2044 32160
rect 2060 32096 2124 32160
rect 2140 32156 2204 32160
rect 2220 32156 2284 32160
rect 2140 32100 2184 32156
rect 2184 32100 2204 32156
rect 2220 32100 2240 32156
rect 2240 32100 2264 32156
rect 2264 32100 2284 32156
rect 2140 32096 2204 32100
rect 2220 32096 2284 32100
rect 7740 32096 7804 32160
rect 7820 32096 7884 32160
rect 7900 32096 7964 32160
rect 7980 32096 8044 32160
rect 8060 32096 8124 32160
rect 8140 32096 8204 32160
rect 8220 32156 8284 32160
rect 8220 32100 8283 32156
rect 8283 32100 8284 32156
rect 8220 32096 8284 32100
rect 13740 32096 13804 32160
rect 13820 32096 13884 32160
rect 13900 32096 13964 32160
rect 13980 32096 14044 32160
rect 14060 32156 14124 32160
rect 14060 32100 14063 32156
rect 14063 32100 14119 32156
rect 14119 32100 14124 32156
rect 14060 32096 14124 32100
rect 14140 32096 14204 32160
rect 14220 32096 14284 32160
rect 19740 32096 19804 32160
rect 19820 32156 19884 32160
rect 19820 32100 19843 32156
rect 19843 32100 19884 32156
rect 19820 32096 19884 32100
rect 19900 32096 19964 32160
rect 19980 32096 20044 32160
rect 20060 32096 20124 32160
rect 20140 32096 20204 32160
rect 20220 32096 20284 32160
rect 25740 32096 25804 32160
rect 25820 32096 25884 32160
rect 25900 32096 25964 32160
rect 25980 32096 26044 32160
rect 26060 32096 26124 32160
rect 26140 32096 26204 32160
rect 26220 32096 26284 32160
rect 31740 32096 31804 32160
rect 31820 32096 31884 32160
rect 31900 32096 31964 32160
rect 31980 32096 32044 32160
rect 32060 32096 32124 32160
rect 32140 32096 32204 32160
rect 32220 32096 32284 32160
rect 37740 32096 37804 32160
rect 37820 32096 37884 32160
rect 37900 32096 37964 32160
rect 37980 32096 38044 32160
rect 38060 32096 38124 32160
rect 38140 32096 38204 32160
rect 38220 32096 38284 32160
rect 43740 32096 43804 32160
rect 43820 32096 43884 32160
rect 43900 32096 43964 32160
rect 43980 32096 44044 32160
rect 44060 32096 44124 32160
rect 44140 32096 44204 32160
rect 44220 32096 44284 32160
rect 49740 32156 49804 32160
rect 49740 32100 49742 32156
rect 49742 32100 49798 32156
rect 49798 32100 49804 32156
rect 49740 32096 49804 32100
rect 49820 32096 49884 32160
rect 49900 32096 49964 32160
rect 49980 32096 50044 32160
rect 50060 32096 50124 32160
rect 50140 32096 50204 32160
rect 50220 32096 50284 32160
rect 55740 32096 55804 32160
rect 55820 32096 55884 32160
rect 55900 32096 55964 32160
rect 55980 32096 56044 32160
rect 56060 32096 56124 32160
rect 56140 32096 56204 32160
rect 56220 32096 56284 32160
rect 61740 32096 61804 32160
rect 61820 32096 61884 32160
rect 61900 32096 61964 32160
rect 61980 32096 62044 32160
rect 62060 32096 62124 32160
rect 62140 32096 62204 32160
rect 62220 32096 62284 32160
rect 67740 32096 67804 32160
rect 67820 32096 67884 32160
rect 67900 32096 67964 32160
rect 67980 32096 68044 32160
rect 68060 32096 68124 32160
rect 68140 32096 68204 32160
rect 68220 32096 68284 32160
rect 73740 32096 73804 32160
rect 73820 32096 73884 32160
rect 73900 32096 73964 32160
rect 73980 32096 74044 32160
rect 74060 32096 74124 32160
rect 74140 32096 74204 32160
rect 74220 32096 74284 32160
rect 1740 32016 1804 32080
rect 1820 32016 1884 32080
rect 1900 32016 1964 32080
rect 1980 32016 2044 32080
rect 2060 32016 2124 32080
rect 2140 32076 2204 32080
rect 2220 32076 2284 32080
rect 2140 32020 2184 32076
rect 2184 32020 2204 32076
rect 2220 32020 2240 32076
rect 2240 32020 2264 32076
rect 2264 32020 2284 32076
rect 2140 32016 2204 32020
rect 2220 32016 2284 32020
rect 7740 32016 7804 32080
rect 7820 32016 7884 32080
rect 7900 32016 7964 32080
rect 7980 32016 8044 32080
rect 8060 32016 8124 32080
rect 8140 32016 8204 32080
rect 8220 32076 8284 32080
rect 8220 32020 8283 32076
rect 8283 32020 8284 32076
rect 8220 32016 8284 32020
rect 13740 32016 13804 32080
rect 13820 32016 13884 32080
rect 13900 32016 13964 32080
rect 13980 32016 14044 32080
rect 14060 32076 14124 32080
rect 14060 32020 14063 32076
rect 14063 32020 14119 32076
rect 14119 32020 14124 32076
rect 14060 32016 14124 32020
rect 14140 32016 14204 32080
rect 14220 32016 14284 32080
rect 19740 32016 19804 32080
rect 19820 32076 19884 32080
rect 19820 32020 19843 32076
rect 19843 32020 19884 32076
rect 19820 32016 19884 32020
rect 19900 32016 19964 32080
rect 19980 32016 20044 32080
rect 20060 32016 20124 32080
rect 20140 32016 20204 32080
rect 20220 32016 20284 32080
rect 25740 32016 25804 32080
rect 25820 32016 25884 32080
rect 25900 32016 25964 32080
rect 25980 32016 26044 32080
rect 26060 32016 26124 32080
rect 26140 32016 26204 32080
rect 26220 32016 26284 32080
rect 31740 32016 31804 32080
rect 31820 32016 31884 32080
rect 31900 32016 31964 32080
rect 31980 32016 32044 32080
rect 32060 32016 32124 32080
rect 32140 32016 32204 32080
rect 32220 32016 32284 32080
rect 37740 32016 37804 32080
rect 37820 32016 37884 32080
rect 37900 32016 37964 32080
rect 37980 32016 38044 32080
rect 38060 32016 38124 32080
rect 38140 32016 38204 32080
rect 38220 32016 38284 32080
rect 43740 32016 43804 32080
rect 43820 32016 43884 32080
rect 43900 32016 43964 32080
rect 43980 32016 44044 32080
rect 44060 32016 44124 32080
rect 44140 32016 44204 32080
rect 44220 32016 44284 32080
rect 49740 32076 49804 32080
rect 49740 32020 49742 32076
rect 49742 32020 49798 32076
rect 49798 32020 49804 32076
rect 49740 32016 49804 32020
rect 49820 32016 49884 32080
rect 49900 32016 49964 32080
rect 49980 32016 50044 32080
rect 50060 32016 50124 32080
rect 50140 32016 50204 32080
rect 50220 32016 50284 32080
rect 55740 32016 55804 32080
rect 55820 32016 55884 32080
rect 55900 32016 55964 32080
rect 55980 32016 56044 32080
rect 56060 32016 56124 32080
rect 56140 32016 56204 32080
rect 56220 32016 56284 32080
rect 61740 32016 61804 32080
rect 61820 32016 61884 32080
rect 61900 32016 61964 32080
rect 61980 32016 62044 32080
rect 62060 32016 62124 32080
rect 62140 32016 62204 32080
rect 62220 32016 62284 32080
rect 67740 32016 67804 32080
rect 67820 32016 67884 32080
rect 67900 32016 67964 32080
rect 67980 32016 68044 32080
rect 68060 32016 68124 32080
rect 68140 32016 68204 32080
rect 68220 32016 68284 32080
rect 73740 32016 73804 32080
rect 73820 32016 73884 32080
rect 73900 32016 73964 32080
rect 73980 32016 74044 32080
rect 74060 32016 74124 32080
rect 74140 32016 74204 32080
rect 74220 32016 74284 32080
rect 1740 31936 1804 32000
rect 1820 31936 1884 32000
rect 1900 31936 1964 32000
rect 1980 31936 2044 32000
rect 2060 31936 2124 32000
rect 2140 31996 2204 32000
rect 2220 31996 2284 32000
rect 2140 31940 2184 31996
rect 2184 31940 2204 31996
rect 2220 31940 2240 31996
rect 2240 31940 2264 31996
rect 2264 31940 2284 31996
rect 2140 31936 2204 31940
rect 2220 31936 2284 31940
rect 7740 31936 7804 32000
rect 7820 31936 7884 32000
rect 7900 31936 7964 32000
rect 7980 31936 8044 32000
rect 8060 31936 8124 32000
rect 8140 31936 8204 32000
rect 8220 31996 8284 32000
rect 8220 31940 8283 31996
rect 8283 31940 8284 31996
rect 8220 31936 8284 31940
rect 13740 31936 13804 32000
rect 13820 31936 13884 32000
rect 13900 31936 13964 32000
rect 13980 31936 14044 32000
rect 14060 31996 14124 32000
rect 14060 31940 14063 31996
rect 14063 31940 14119 31996
rect 14119 31940 14124 31996
rect 14060 31936 14124 31940
rect 14140 31936 14204 32000
rect 14220 31936 14284 32000
rect 19740 31936 19804 32000
rect 19820 31996 19884 32000
rect 19820 31940 19843 31996
rect 19843 31940 19884 31996
rect 19820 31936 19884 31940
rect 19900 31936 19964 32000
rect 19980 31936 20044 32000
rect 20060 31936 20124 32000
rect 20140 31936 20204 32000
rect 20220 31936 20284 32000
rect 25740 31936 25804 32000
rect 25820 31936 25884 32000
rect 25900 31936 25964 32000
rect 25980 31936 26044 32000
rect 26060 31936 26124 32000
rect 26140 31936 26204 32000
rect 26220 31936 26284 32000
rect 31740 31936 31804 32000
rect 31820 31936 31884 32000
rect 31900 31936 31964 32000
rect 31980 31936 32044 32000
rect 32060 31936 32124 32000
rect 32140 31936 32204 32000
rect 32220 31936 32284 32000
rect 37740 31936 37804 32000
rect 37820 31936 37884 32000
rect 37900 31936 37964 32000
rect 37980 31936 38044 32000
rect 38060 31936 38124 32000
rect 38140 31936 38204 32000
rect 38220 31936 38284 32000
rect 43740 31936 43804 32000
rect 43820 31936 43884 32000
rect 43900 31936 43964 32000
rect 43980 31936 44044 32000
rect 44060 31936 44124 32000
rect 44140 31936 44204 32000
rect 44220 31936 44284 32000
rect 49740 31996 49804 32000
rect 49740 31940 49742 31996
rect 49742 31940 49798 31996
rect 49798 31940 49804 31996
rect 49740 31936 49804 31940
rect 49820 31936 49884 32000
rect 49900 31936 49964 32000
rect 49980 31936 50044 32000
rect 50060 31936 50124 32000
rect 50140 31936 50204 32000
rect 50220 31936 50284 32000
rect 55740 31936 55804 32000
rect 55820 31936 55884 32000
rect 55900 31936 55964 32000
rect 55980 31936 56044 32000
rect 56060 31936 56124 32000
rect 56140 31936 56204 32000
rect 56220 31936 56284 32000
rect 61740 31936 61804 32000
rect 61820 31936 61884 32000
rect 61900 31936 61964 32000
rect 61980 31936 62044 32000
rect 62060 31936 62124 32000
rect 62140 31936 62204 32000
rect 62220 31936 62284 32000
rect 67740 31936 67804 32000
rect 67820 31936 67884 32000
rect 67900 31936 67964 32000
rect 67980 31936 68044 32000
rect 68060 31936 68124 32000
rect 68140 31936 68204 32000
rect 68220 31936 68284 32000
rect 73740 31936 73804 32000
rect 73820 31936 73884 32000
rect 73900 31936 73964 32000
rect 73980 31936 74044 32000
rect 74060 31936 74124 32000
rect 74140 31936 74204 32000
rect 74220 31936 74284 32000
rect 4740 24528 4804 24592
rect 4820 24528 4884 24592
rect 4900 24528 4964 24592
rect 4980 24528 5044 24592
rect 5060 24528 5124 24592
rect 5140 24528 5204 24592
rect 5220 24528 5284 24592
rect 10740 24528 10804 24592
rect 10820 24528 10884 24592
rect 10900 24528 10964 24592
rect 10980 24528 11044 24592
rect 11060 24528 11124 24592
rect 11140 24528 11204 24592
rect 11220 24528 11284 24592
rect 16740 24528 16804 24592
rect 16820 24528 16884 24592
rect 16900 24528 16964 24592
rect 16980 24528 17044 24592
rect 17060 24588 17124 24592
rect 17140 24588 17204 24592
rect 17060 24532 17100 24588
rect 17100 24532 17124 24588
rect 17140 24532 17156 24588
rect 17156 24532 17204 24588
rect 17060 24528 17124 24532
rect 17140 24528 17204 24532
rect 17220 24528 17284 24592
rect 22740 24528 22804 24592
rect 22820 24588 22884 24592
rect 22900 24588 22964 24592
rect 22820 24532 22880 24588
rect 22880 24532 22884 24588
rect 22900 24532 22936 24588
rect 22936 24532 22964 24588
rect 22820 24528 22884 24532
rect 22900 24528 22964 24532
rect 22980 24528 23044 24592
rect 23060 24528 23124 24592
rect 23140 24528 23204 24592
rect 23220 24528 23284 24592
rect 28740 24528 28804 24592
rect 28820 24528 28884 24592
rect 28900 24528 28964 24592
rect 28980 24528 29044 24592
rect 29060 24528 29124 24592
rect 29140 24528 29204 24592
rect 29220 24528 29284 24592
rect 34740 24528 34804 24592
rect 34820 24528 34884 24592
rect 34900 24528 34964 24592
rect 34980 24528 35044 24592
rect 35060 24528 35124 24592
rect 35140 24528 35204 24592
rect 35220 24528 35284 24592
rect 40740 24528 40804 24592
rect 40820 24528 40884 24592
rect 40900 24528 40964 24592
rect 40980 24528 41044 24592
rect 41060 24528 41124 24592
rect 41140 24528 41204 24592
rect 41220 24528 41284 24592
rect 46740 24528 46804 24592
rect 46820 24528 46884 24592
rect 46900 24528 46964 24592
rect 46980 24528 47044 24592
rect 47060 24528 47124 24592
rect 47140 24528 47204 24592
rect 47220 24528 47284 24592
rect 52740 24528 52804 24592
rect 52820 24528 52884 24592
rect 52900 24528 52964 24592
rect 52980 24528 53044 24592
rect 53060 24528 53124 24592
rect 53140 24528 53204 24592
rect 53220 24528 53284 24592
rect 58740 24528 58804 24592
rect 58820 24528 58884 24592
rect 58900 24528 58964 24592
rect 58980 24528 59044 24592
rect 59060 24588 59124 24592
rect 59060 24532 59104 24588
rect 59104 24532 59124 24588
rect 59060 24528 59124 24532
rect 59140 24528 59204 24592
rect 59220 24528 59284 24592
rect 64740 24528 64804 24592
rect 64820 24528 64884 24592
rect 64900 24528 64964 24592
rect 64980 24528 65044 24592
rect 65060 24528 65124 24592
rect 65140 24528 65204 24592
rect 65220 24528 65284 24592
rect 70740 24528 70804 24592
rect 70820 24528 70884 24592
rect 70900 24528 70964 24592
rect 70980 24528 71044 24592
rect 71060 24528 71124 24592
rect 71140 24528 71204 24592
rect 71220 24528 71284 24592
rect 4740 24448 4804 24512
rect 4820 24448 4884 24512
rect 4900 24448 4964 24512
rect 4980 24448 5044 24512
rect 5060 24448 5124 24512
rect 5140 24448 5204 24512
rect 5220 24448 5284 24512
rect 10740 24448 10804 24512
rect 10820 24448 10884 24512
rect 10900 24448 10964 24512
rect 10980 24448 11044 24512
rect 11060 24448 11124 24512
rect 11140 24448 11204 24512
rect 11220 24448 11284 24512
rect 16740 24448 16804 24512
rect 16820 24448 16884 24512
rect 16900 24448 16964 24512
rect 16980 24448 17044 24512
rect 17060 24508 17124 24512
rect 17140 24508 17204 24512
rect 17060 24452 17100 24508
rect 17100 24452 17124 24508
rect 17140 24452 17156 24508
rect 17156 24452 17204 24508
rect 17060 24448 17124 24452
rect 17140 24448 17204 24452
rect 17220 24448 17284 24512
rect 22740 24448 22804 24512
rect 22820 24508 22884 24512
rect 22900 24508 22964 24512
rect 22820 24452 22880 24508
rect 22880 24452 22884 24508
rect 22900 24452 22936 24508
rect 22936 24452 22964 24508
rect 22820 24448 22884 24452
rect 22900 24448 22964 24452
rect 22980 24448 23044 24512
rect 23060 24448 23124 24512
rect 23140 24448 23204 24512
rect 23220 24448 23284 24512
rect 28740 24448 28804 24512
rect 28820 24448 28884 24512
rect 28900 24448 28964 24512
rect 28980 24448 29044 24512
rect 29060 24448 29124 24512
rect 29140 24448 29204 24512
rect 29220 24448 29284 24512
rect 34740 24448 34804 24512
rect 34820 24448 34884 24512
rect 34900 24448 34964 24512
rect 34980 24448 35044 24512
rect 35060 24448 35124 24512
rect 35140 24448 35204 24512
rect 35220 24448 35284 24512
rect 40740 24448 40804 24512
rect 40820 24448 40884 24512
rect 40900 24448 40964 24512
rect 40980 24448 41044 24512
rect 41060 24448 41124 24512
rect 41140 24448 41204 24512
rect 41220 24448 41284 24512
rect 46740 24448 46804 24512
rect 46820 24448 46884 24512
rect 46900 24448 46964 24512
rect 46980 24448 47044 24512
rect 47060 24448 47124 24512
rect 47140 24448 47204 24512
rect 47220 24448 47284 24512
rect 52740 24448 52804 24512
rect 52820 24448 52884 24512
rect 52900 24448 52964 24512
rect 52980 24448 53044 24512
rect 53060 24448 53124 24512
rect 53140 24448 53204 24512
rect 53220 24448 53284 24512
rect 58740 24448 58804 24512
rect 58820 24448 58884 24512
rect 58900 24448 58964 24512
rect 58980 24448 59044 24512
rect 59060 24508 59124 24512
rect 59060 24452 59104 24508
rect 59104 24452 59124 24508
rect 59060 24448 59124 24452
rect 59140 24448 59204 24512
rect 59220 24448 59284 24512
rect 64740 24448 64804 24512
rect 64820 24448 64884 24512
rect 64900 24448 64964 24512
rect 64980 24448 65044 24512
rect 65060 24448 65124 24512
rect 65140 24448 65204 24512
rect 65220 24448 65284 24512
rect 70740 24448 70804 24512
rect 70820 24448 70884 24512
rect 70900 24448 70964 24512
rect 70980 24448 71044 24512
rect 71060 24448 71124 24512
rect 71140 24448 71204 24512
rect 71220 24448 71284 24512
rect 4740 24368 4804 24432
rect 4820 24368 4884 24432
rect 4900 24368 4964 24432
rect 4980 24368 5044 24432
rect 5060 24368 5124 24432
rect 5140 24368 5204 24432
rect 5220 24368 5284 24432
rect 10740 24368 10804 24432
rect 10820 24368 10884 24432
rect 10900 24368 10964 24432
rect 10980 24368 11044 24432
rect 11060 24368 11124 24432
rect 11140 24368 11204 24432
rect 11220 24368 11284 24432
rect 16740 24368 16804 24432
rect 16820 24368 16884 24432
rect 16900 24368 16964 24432
rect 16980 24368 17044 24432
rect 17060 24428 17124 24432
rect 17140 24428 17204 24432
rect 17060 24372 17100 24428
rect 17100 24372 17124 24428
rect 17140 24372 17156 24428
rect 17156 24372 17204 24428
rect 17060 24368 17124 24372
rect 17140 24368 17204 24372
rect 17220 24368 17284 24432
rect 22740 24368 22804 24432
rect 22820 24428 22884 24432
rect 22900 24428 22964 24432
rect 22820 24372 22880 24428
rect 22880 24372 22884 24428
rect 22900 24372 22936 24428
rect 22936 24372 22964 24428
rect 22820 24368 22884 24372
rect 22900 24368 22964 24372
rect 22980 24368 23044 24432
rect 23060 24368 23124 24432
rect 23140 24368 23204 24432
rect 23220 24368 23284 24432
rect 28740 24368 28804 24432
rect 28820 24368 28884 24432
rect 28900 24368 28964 24432
rect 28980 24368 29044 24432
rect 29060 24368 29124 24432
rect 29140 24368 29204 24432
rect 29220 24368 29284 24432
rect 34740 24368 34804 24432
rect 34820 24368 34884 24432
rect 34900 24368 34964 24432
rect 34980 24368 35044 24432
rect 35060 24368 35124 24432
rect 35140 24368 35204 24432
rect 35220 24368 35284 24432
rect 40740 24368 40804 24432
rect 40820 24368 40884 24432
rect 40900 24368 40964 24432
rect 40980 24368 41044 24432
rect 41060 24368 41124 24432
rect 41140 24368 41204 24432
rect 41220 24368 41284 24432
rect 46740 24368 46804 24432
rect 46820 24368 46884 24432
rect 46900 24368 46964 24432
rect 46980 24368 47044 24432
rect 47060 24368 47124 24432
rect 47140 24368 47204 24432
rect 47220 24368 47284 24432
rect 52740 24368 52804 24432
rect 52820 24368 52884 24432
rect 52900 24368 52964 24432
rect 52980 24368 53044 24432
rect 53060 24368 53124 24432
rect 53140 24368 53204 24432
rect 53220 24368 53284 24432
rect 58740 24368 58804 24432
rect 58820 24368 58884 24432
rect 58900 24368 58964 24432
rect 58980 24368 59044 24432
rect 59060 24428 59124 24432
rect 59060 24372 59104 24428
rect 59104 24372 59124 24428
rect 59060 24368 59124 24372
rect 59140 24368 59204 24432
rect 59220 24368 59284 24432
rect 64740 24368 64804 24432
rect 64820 24368 64884 24432
rect 64900 24368 64964 24432
rect 64980 24368 65044 24432
rect 65060 24368 65124 24432
rect 65140 24368 65204 24432
rect 65220 24368 65284 24432
rect 70740 24368 70804 24432
rect 70820 24368 70884 24432
rect 70900 24368 70964 24432
rect 70980 24368 71044 24432
rect 71060 24368 71124 24432
rect 71140 24368 71204 24432
rect 71220 24368 71284 24432
rect 4740 24288 4804 24352
rect 4820 24288 4884 24352
rect 4900 24288 4964 24352
rect 4980 24288 5044 24352
rect 5060 24288 5124 24352
rect 5140 24288 5204 24352
rect 5220 24288 5284 24352
rect 10740 24288 10804 24352
rect 10820 24288 10884 24352
rect 10900 24288 10964 24352
rect 10980 24288 11044 24352
rect 11060 24288 11124 24352
rect 11140 24288 11204 24352
rect 11220 24288 11284 24352
rect 16740 24288 16804 24352
rect 16820 24288 16884 24352
rect 16900 24288 16964 24352
rect 16980 24288 17044 24352
rect 17060 24348 17124 24352
rect 17140 24348 17204 24352
rect 17060 24292 17100 24348
rect 17100 24292 17124 24348
rect 17140 24292 17156 24348
rect 17156 24292 17204 24348
rect 17060 24288 17124 24292
rect 17140 24288 17204 24292
rect 17220 24288 17284 24352
rect 22740 24288 22804 24352
rect 22820 24348 22884 24352
rect 22900 24348 22964 24352
rect 22820 24292 22880 24348
rect 22880 24292 22884 24348
rect 22900 24292 22936 24348
rect 22936 24292 22964 24348
rect 22820 24288 22884 24292
rect 22900 24288 22964 24292
rect 22980 24288 23044 24352
rect 23060 24288 23124 24352
rect 23140 24288 23204 24352
rect 23220 24288 23284 24352
rect 28740 24288 28804 24352
rect 28820 24288 28884 24352
rect 28900 24288 28964 24352
rect 28980 24288 29044 24352
rect 29060 24288 29124 24352
rect 29140 24288 29204 24352
rect 29220 24288 29284 24352
rect 34740 24288 34804 24352
rect 34820 24288 34884 24352
rect 34900 24288 34964 24352
rect 34980 24288 35044 24352
rect 35060 24288 35124 24352
rect 35140 24288 35204 24352
rect 35220 24288 35284 24352
rect 40740 24288 40804 24352
rect 40820 24288 40884 24352
rect 40900 24288 40964 24352
rect 40980 24288 41044 24352
rect 41060 24288 41124 24352
rect 41140 24288 41204 24352
rect 41220 24288 41284 24352
rect 46740 24288 46804 24352
rect 46820 24288 46884 24352
rect 46900 24288 46964 24352
rect 46980 24288 47044 24352
rect 47060 24288 47124 24352
rect 47140 24288 47204 24352
rect 47220 24288 47284 24352
rect 52740 24288 52804 24352
rect 52820 24288 52884 24352
rect 52900 24288 52964 24352
rect 52980 24288 53044 24352
rect 53060 24288 53124 24352
rect 53140 24288 53204 24352
rect 53220 24288 53284 24352
rect 58740 24288 58804 24352
rect 58820 24288 58884 24352
rect 58900 24288 58964 24352
rect 58980 24288 59044 24352
rect 59060 24348 59124 24352
rect 59060 24292 59104 24348
rect 59104 24292 59124 24348
rect 59060 24288 59124 24292
rect 59140 24288 59204 24352
rect 59220 24288 59284 24352
rect 64740 24288 64804 24352
rect 64820 24288 64884 24352
rect 64900 24288 64964 24352
rect 64980 24288 65044 24352
rect 65060 24288 65124 24352
rect 65140 24288 65204 24352
rect 65220 24288 65284 24352
rect 70740 24288 70804 24352
rect 70820 24288 70884 24352
rect 70900 24288 70964 24352
rect 70980 24288 71044 24352
rect 71060 24288 71124 24352
rect 71140 24288 71204 24352
rect 71220 24288 71284 24352
rect 66300 23488 66364 23492
rect 66300 23432 66350 23488
rect 66350 23432 66364 23488
rect 66300 23428 66364 23432
rect 66484 23488 66548 23492
rect 66484 23432 66534 23488
rect 66534 23432 66548 23488
rect 66484 23428 66548 23432
rect 1740 22176 1804 22240
rect 1820 22176 1884 22240
rect 1900 22176 1964 22240
rect 1980 22176 2044 22240
rect 2060 22176 2124 22240
rect 2140 22236 2204 22240
rect 2220 22236 2284 22240
rect 2140 22180 2184 22236
rect 2184 22180 2204 22236
rect 2220 22180 2240 22236
rect 2240 22180 2264 22236
rect 2264 22180 2284 22236
rect 2140 22176 2204 22180
rect 2220 22176 2284 22180
rect 7740 22176 7804 22240
rect 7820 22176 7884 22240
rect 7900 22176 7964 22240
rect 7980 22176 8044 22240
rect 8060 22176 8124 22240
rect 8140 22176 8204 22240
rect 8220 22236 8284 22240
rect 8220 22180 8283 22236
rect 8283 22180 8284 22236
rect 8220 22176 8284 22180
rect 13740 22176 13804 22240
rect 13820 22176 13884 22240
rect 13900 22176 13964 22240
rect 13980 22176 14044 22240
rect 14060 22236 14124 22240
rect 14060 22180 14063 22236
rect 14063 22180 14119 22236
rect 14119 22180 14124 22236
rect 14060 22176 14124 22180
rect 14140 22176 14204 22240
rect 14220 22176 14284 22240
rect 19740 22176 19804 22240
rect 19820 22236 19884 22240
rect 19820 22180 19843 22236
rect 19843 22180 19884 22236
rect 19820 22176 19884 22180
rect 19900 22176 19964 22240
rect 19980 22176 20044 22240
rect 20060 22176 20124 22240
rect 20140 22176 20204 22240
rect 20220 22176 20284 22240
rect 25740 22176 25804 22240
rect 25820 22176 25884 22240
rect 25900 22176 25964 22240
rect 25980 22176 26044 22240
rect 26060 22176 26124 22240
rect 26140 22176 26204 22240
rect 26220 22176 26284 22240
rect 31740 22176 31804 22240
rect 31820 22176 31884 22240
rect 31900 22176 31964 22240
rect 31980 22176 32044 22240
rect 32060 22176 32124 22240
rect 32140 22176 32204 22240
rect 32220 22176 32284 22240
rect 37740 22176 37804 22240
rect 37820 22176 37884 22240
rect 37900 22176 37964 22240
rect 37980 22176 38044 22240
rect 38060 22176 38124 22240
rect 38140 22176 38204 22240
rect 38220 22176 38284 22240
rect 43740 22176 43804 22240
rect 43820 22176 43884 22240
rect 43900 22176 43964 22240
rect 43980 22176 44044 22240
rect 44060 22176 44124 22240
rect 44140 22176 44204 22240
rect 44220 22176 44284 22240
rect 49740 22236 49804 22240
rect 49740 22180 49742 22236
rect 49742 22180 49798 22236
rect 49798 22180 49804 22236
rect 49740 22176 49804 22180
rect 49820 22176 49884 22240
rect 49900 22176 49964 22240
rect 49980 22176 50044 22240
rect 50060 22176 50124 22240
rect 50140 22176 50204 22240
rect 50220 22176 50284 22240
rect 55740 22176 55804 22240
rect 55820 22176 55884 22240
rect 55900 22176 55964 22240
rect 55980 22176 56044 22240
rect 56060 22176 56124 22240
rect 56140 22176 56204 22240
rect 56220 22176 56284 22240
rect 61740 22176 61804 22240
rect 61820 22176 61884 22240
rect 61900 22176 61964 22240
rect 61980 22176 62044 22240
rect 62060 22176 62124 22240
rect 62140 22176 62204 22240
rect 62220 22176 62284 22240
rect 67740 22176 67804 22240
rect 67820 22176 67884 22240
rect 67900 22176 67964 22240
rect 67980 22176 68044 22240
rect 68060 22176 68124 22240
rect 68140 22176 68204 22240
rect 68220 22176 68284 22240
rect 73740 22176 73804 22240
rect 73820 22176 73884 22240
rect 73900 22176 73964 22240
rect 73980 22176 74044 22240
rect 74060 22176 74124 22240
rect 74140 22176 74204 22240
rect 74220 22176 74284 22240
rect 1740 22096 1804 22160
rect 1820 22096 1884 22160
rect 1900 22096 1964 22160
rect 1980 22096 2044 22160
rect 2060 22096 2124 22160
rect 2140 22156 2204 22160
rect 2220 22156 2284 22160
rect 2140 22100 2184 22156
rect 2184 22100 2204 22156
rect 2220 22100 2240 22156
rect 2240 22100 2264 22156
rect 2264 22100 2284 22156
rect 2140 22096 2204 22100
rect 2220 22096 2284 22100
rect 7740 22096 7804 22160
rect 7820 22096 7884 22160
rect 7900 22096 7964 22160
rect 7980 22096 8044 22160
rect 8060 22096 8124 22160
rect 8140 22096 8204 22160
rect 8220 22156 8284 22160
rect 8220 22100 8283 22156
rect 8283 22100 8284 22156
rect 8220 22096 8284 22100
rect 13740 22096 13804 22160
rect 13820 22096 13884 22160
rect 13900 22096 13964 22160
rect 13980 22096 14044 22160
rect 14060 22156 14124 22160
rect 14060 22100 14063 22156
rect 14063 22100 14119 22156
rect 14119 22100 14124 22156
rect 14060 22096 14124 22100
rect 14140 22096 14204 22160
rect 14220 22096 14284 22160
rect 19740 22096 19804 22160
rect 19820 22156 19884 22160
rect 19820 22100 19843 22156
rect 19843 22100 19884 22156
rect 19820 22096 19884 22100
rect 19900 22096 19964 22160
rect 19980 22096 20044 22160
rect 20060 22096 20124 22160
rect 20140 22096 20204 22160
rect 20220 22096 20284 22160
rect 25740 22096 25804 22160
rect 25820 22096 25884 22160
rect 25900 22096 25964 22160
rect 25980 22096 26044 22160
rect 26060 22096 26124 22160
rect 26140 22096 26204 22160
rect 26220 22096 26284 22160
rect 31740 22096 31804 22160
rect 31820 22096 31884 22160
rect 31900 22096 31964 22160
rect 31980 22096 32044 22160
rect 32060 22096 32124 22160
rect 32140 22096 32204 22160
rect 32220 22096 32284 22160
rect 37740 22096 37804 22160
rect 37820 22096 37884 22160
rect 37900 22096 37964 22160
rect 37980 22096 38044 22160
rect 38060 22096 38124 22160
rect 38140 22096 38204 22160
rect 38220 22096 38284 22160
rect 43740 22096 43804 22160
rect 43820 22096 43884 22160
rect 43900 22096 43964 22160
rect 43980 22096 44044 22160
rect 44060 22096 44124 22160
rect 44140 22096 44204 22160
rect 44220 22096 44284 22160
rect 49740 22156 49804 22160
rect 49740 22100 49742 22156
rect 49742 22100 49798 22156
rect 49798 22100 49804 22156
rect 49740 22096 49804 22100
rect 49820 22096 49884 22160
rect 49900 22096 49964 22160
rect 49980 22096 50044 22160
rect 50060 22096 50124 22160
rect 50140 22096 50204 22160
rect 50220 22096 50284 22160
rect 55740 22096 55804 22160
rect 55820 22096 55884 22160
rect 55900 22096 55964 22160
rect 55980 22096 56044 22160
rect 56060 22096 56124 22160
rect 56140 22096 56204 22160
rect 56220 22096 56284 22160
rect 61740 22096 61804 22160
rect 61820 22096 61884 22160
rect 61900 22096 61964 22160
rect 61980 22096 62044 22160
rect 62060 22096 62124 22160
rect 62140 22096 62204 22160
rect 62220 22096 62284 22160
rect 67740 22096 67804 22160
rect 67820 22096 67884 22160
rect 67900 22096 67964 22160
rect 67980 22096 68044 22160
rect 68060 22096 68124 22160
rect 68140 22096 68204 22160
rect 68220 22096 68284 22160
rect 73740 22096 73804 22160
rect 73820 22096 73884 22160
rect 73900 22096 73964 22160
rect 73980 22096 74044 22160
rect 74060 22096 74124 22160
rect 74140 22096 74204 22160
rect 74220 22096 74284 22160
rect 1740 22016 1804 22080
rect 1820 22016 1884 22080
rect 1900 22016 1964 22080
rect 1980 22016 2044 22080
rect 2060 22016 2124 22080
rect 2140 22076 2204 22080
rect 2220 22076 2284 22080
rect 2140 22020 2184 22076
rect 2184 22020 2204 22076
rect 2220 22020 2240 22076
rect 2240 22020 2264 22076
rect 2264 22020 2284 22076
rect 2140 22016 2204 22020
rect 2220 22016 2284 22020
rect 7740 22016 7804 22080
rect 7820 22016 7884 22080
rect 7900 22016 7964 22080
rect 7980 22016 8044 22080
rect 8060 22016 8124 22080
rect 8140 22016 8204 22080
rect 8220 22076 8284 22080
rect 8220 22020 8283 22076
rect 8283 22020 8284 22076
rect 8220 22016 8284 22020
rect 13740 22016 13804 22080
rect 13820 22016 13884 22080
rect 13900 22016 13964 22080
rect 13980 22016 14044 22080
rect 14060 22076 14124 22080
rect 14060 22020 14063 22076
rect 14063 22020 14119 22076
rect 14119 22020 14124 22076
rect 14060 22016 14124 22020
rect 14140 22016 14204 22080
rect 14220 22016 14284 22080
rect 19740 22016 19804 22080
rect 19820 22076 19884 22080
rect 19820 22020 19843 22076
rect 19843 22020 19884 22076
rect 19820 22016 19884 22020
rect 19900 22016 19964 22080
rect 19980 22016 20044 22080
rect 20060 22016 20124 22080
rect 20140 22016 20204 22080
rect 20220 22016 20284 22080
rect 25740 22016 25804 22080
rect 25820 22016 25884 22080
rect 25900 22016 25964 22080
rect 25980 22016 26044 22080
rect 26060 22016 26124 22080
rect 26140 22016 26204 22080
rect 26220 22016 26284 22080
rect 31740 22016 31804 22080
rect 31820 22016 31884 22080
rect 31900 22016 31964 22080
rect 31980 22016 32044 22080
rect 32060 22016 32124 22080
rect 32140 22016 32204 22080
rect 32220 22016 32284 22080
rect 37740 22016 37804 22080
rect 37820 22016 37884 22080
rect 37900 22016 37964 22080
rect 37980 22016 38044 22080
rect 38060 22016 38124 22080
rect 38140 22016 38204 22080
rect 38220 22016 38284 22080
rect 43740 22016 43804 22080
rect 43820 22016 43884 22080
rect 43900 22016 43964 22080
rect 43980 22016 44044 22080
rect 44060 22016 44124 22080
rect 44140 22016 44204 22080
rect 44220 22016 44284 22080
rect 49740 22076 49804 22080
rect 49740 22020 49742 22076
rect 49742 22020 49798 22076
rect 49798 22020 49804 22076
rect 49740 22016 49804 22020
rect 49820 22016 49884 22080
rect 49900 22016 49964 22080
rect 49980 22016 50044 22080
rect 50060 22016 50124 22080
rect 50140 22016 50204 22080
rect 50220 22016 50284 22080
rect 55740 22016 55804 22080
rect 55820 22016 55884 22080
rect 55900 22016 55964 22080
rect 55980 22016 56044 22080
rect 56060 22016 56124 22080
rect 56140 22016 56204 22080
rect 56220 22016 56284 22080
rect 61740 22016 61804 22080
rect 61820 22016 61884 22080
rect 61900 22016 61964 22080
rect 61980 22016 62044 22080
rect 62060 22016 62124 22080
rect 62140 22016 62204 22080
rect 62220 22016 62284 22080
rect 67740 22016 67804 22080
rect 67820 22016 67884 22080
rect 67900 22016 67964 22080
rect 67980 22016 68044 22080
rect 68060 22016 68124 22080
rect 68140 22016 68204 22080
rect 68220 22016 68284 22080
rect 73740 22016 73804 22080
rect 73820 22016 73884 22080
rect 73900 22016 73964 22080
rect 73980 22016 74044 22080
rect 74060 22016 74124 22080
rect 74140 22016 74204 22080
rect 74220 22016 74284 22080
rect 1740 21936 1804 22000
rect 1820 21936 1884 22000
rect 1900 21936 1964 22000
rect 1980 21936 2044 22000
rect 2060 21936 2124 22000
rect 2140 21996 2204 22000
rect 2220 21996 2284 22000
rect 2140 21940 2184 21996
rect 2184 21940 2204 21996
rect 2220 21940 2240 21996
rect 2240 21940 2264 21996
rect 2264 21940 2284 21996
rect 2140 21936 2204 21940
rect 2220 21936 2284 21940
rect 7740 21936 7804 22000
rect 7820 21936 7884 22000
rect 7900 21936 7964 22000
rect 7980 21936 8044 22000
rect 8060 21936 8124 22000
rect 8140 21936 8204 22000
rect 8220 21996 8284 22000
rect 8220 21940 8283 21996
rect 8283 21940 8284 21996
rect 8220 21936 8284 21940
rect 13740 21936 13804 22000
rect 13820 21936 13884 22000
rect 13900 21936 13964 22000
rect 13980 21936 14044 22000
rect 14060 21996 14124 22000
rect 14060 21940 14063 21996
rect 14063 21940 14119 21996
rect 14119 21940 14124 21996
rect 14060 21936 14124 21940
rect 14140 21936 14204 22000
rect 14220 21936 14284 22000
rect 19740 21936 19804 22000
rect 19820 21996 19884 22000
rect 19820 21940 19843 21996
rect 19843 21940 19884 21996
rect 19820 21936 19884 21940
rect 19900 21936 19964 22000
rect 19980 21936 20044 22000
rect 20060 21936 20124 22000
rect 20140 21936 20204 22000
rect 20220 21936 20284 22000
rect 25740 21936 25804 22000
rect 25820 21936 25884 22000
rect 25900 21936 25964 22000
rect 25980 21936 26044 22000
rect 26060 21936 26124 22000
rect 26140 21936 26204 22000
rect 26220 21936 26284 22000
rect 31740 21936 31804 22000
rect 31820 21936 31884 22000
rect 31900 21936 31964 22000
rect 31980 21936 32044 22000
rect 32060 21936 32124 22000
rect 32140 21936 32204 22000
rect 32220 21936 32284 22000
rect 37740 21936 37804 22000
rect 37820 21936 37884 22000
rect 37900 21936 37964 22000
rect 37980 21936 38044 22000
rect 38060 21936 38124 22000
rect 38140 21936 38204 22000
rect 38220 21936 38284 22000
rect 43740 21936 43804 22000
rect 43820 21936 43884 22000
rect 43900 21936 43964 22000
rect 43980 21936 44044 22000
rect 44060 21936 44124 22000
rect 44140 21936 44204 22000
rect 44220 21936 44284 22000
rect 49740 21996 49804 22000
rect 49740 21940 49742 21996
rect 49742 21940 49798 21996
rect 49798 21940 49804 21996
rect 49740 21936 49804 21940
rect 49820 21936 49884 22000
rect 49900 21936 49964 22000
rect 49980 21936 50044 22000
rect 50060 21936 50124 22000
rect 50140 21936 50204 22000
rect 50220 21936 50284 22000
rect 55740 21936 55804 22000
rect 55820 21936 55884 22000
rect 55900 21936 55964 22000
rect 55980 21936 56044 22000
rect 56060 21936 56124 22000
rect 56140 21936 56204 22000
rect 56220 21936 56284 22000
rect 61740 21936 61804 22000
rect 61820 21936 61884 22000
rect 61900 21936 61964 22000
rect 61980 21936 62044 22000
rect 62060 21936 62124 22000
rect 62140 21936 62204 22000
rect 62220 21936 62284 22000
rect 67740 21936 67804 22000
rect 67820 21936 67884 22000
rect 67900 21936 67964 22000
rect 67980 21936 68044 22000
rect 68060 21936 68124 22000
rect 68140 21936 68204 22000
rect 68220 21936 68284 22000
rect 73740 21936 73804 22000
rect 73820 21936 73884 22000
rect 73900 21936 73964 22000
rect 73980 21936 74044 22000
rect 74060 21936 74124 22000
rect 74140 21936 74204 22000
rect 74220 21936 74284 22000
rect 66668 19076 66732 19140
rect 62988 17852 63052 17916
rect 4740 14528 4804 14592
rect 4820 14528 4884 14592
rect 4900 14528 4964 14592
rect 4980 14528 5044 14592
rect 5060 14528 5124 14592
rect 5140 14528 5204 14592
rect 5220 14528 5284 14592
rect 10740 14528 10804 14592
rect 10820 14528 10884 14592
rect 10900 14528 10964 14592
rect 10980 14528 11044 14592
rect 11060 14528 11124 14592
rect 11140 14528 11204 14592
rect 11220 14528 11284 14592
rect 16740 14528 16804 14592
rect 16820 14528 16884 14592
rect 16900 14528 16964 14592
rect 16980 14528 17044 14592
rect 17060 14588 17124 14592
rect 17140 14588 17204 14592
rect 17060 14532 17100 14588
rect 17100 14532 17124 14588
rect 17140 14532 17156 14588
rect 17156 14532 17204 14588
rect 17060 14528 17124 14532
rect 17140 14528 17204 14532
rect 17220 14528 17284 14592
rect 22740 14528 22804 14592
rect 22820 14588 22884 14592
rect 22900 14588 22964 14592
rect 22820 14532 22880 14588
rect 22880 14532 22884 14588
rect 22900 14532 22936 14588
rect 22936 14532 22964 14588
rect 22820 14528 22884 14532
rect 22900 14528 22964 14532
rect 22980 14528 23044 14592
rect 23060 14528 23124 14592
rect 23140 14528 23204 14592
rect 23220 14528 23284 14592
rect 28740 14528 28804 14592
rect 28820 14528 28884 14592
rect 28900 14528 28964 14592
rect 28980 14528 29044 14592
rect 29060 14528 29124 14592
rect 29140 14528 29204 14592
rect 29220 14528 29284 14592
rect 34740 14528 34804 14592
rect 34820 14528 34884 14592
rect 34900 14528 34964 14592
rect 34980 14528 35044 14592
rect 35060 14528 35124 14592
rect 35140 14528 35204 14592
rect 35220 14528 35284 14592
rect 40740 14528 40804 14592
rect 40820 14528 40884 14592
rect 40900 14528 40964 14592
rect 40980 14528 41044 14592
rect 41060 14528 41124 14592
rect 41140 14528 41204 14592
rect 41220 14528 41284 14592
rect 46740 14528 46804 14592
rect 46820 14528 46884 14592
rect 46900 14528 46964 14592
rect 46980 14528 47044 14592
rect 47060 14528 47124 14592
rect 47140 14528 47204 14592
rect 47220 14528 47284 14592
rect 52740 14528 52804 14592
rect 52820 14528 52884 14592
rect 52900 14528 52964 14592
rect 52980 14528 53044 14592
rect 53060 14528 53124 14592
rect 53140 14528 53204 14592
rect 53220 14528 53284 14592
rect 58740 14528 58804 14592
rect 58820 14528 58884 14592
rect 58900 14528 58964 14592
rect 58980 14528 59044 14592
rect 59060 14588 59124 14592
rect 59060 14532 59104 14588
rect 59104 14532 59124 14588
rect 59060 14528 59124 14532
rect 59140 14528 59204 14592
rect 59220 14528 59284 14592
rect 64740 14528 64804 14592
rect 64820 14528 64884 14592
rect 64900 14528 64964 14592
rect 64980 14528 65044 14592
rect 65060 14528 65124 14592
rect 65140 14528 65204 14592
rect 65220 14528 65284 14592
rect 70740 14528 70804 14592
rect 70820 14528 70884 14592
rect 70900 14528 70964 14592
rect 70980 14528 71044 14592
rect 71060 14528 71124 14592
rect 71140 14528 71204 14592
rect 71220 14528 71284 14592
rect 4740 14448 4804 14512
rect 4820 14448 4884 14512
rect 4900 14448 4964 14512
rect 4980 14448 5044 14512
rect 5060 14448 5124 14512
rect 5140 14448 5204 14512
rect 5220 14448 5284 14512
rect 10740 14448 10804 14512
rect 10820 14448 10884 14512
rect 10900 14448 10964 14512
rect 10980 14448 11044 14512
rect 11060 14448 11124 14512
rect 11140 14448 11204 14512
rect 11220 14448 11284 14512
rect 16740 14448 16804 14512
rect 16820 14448 16884 14512
rect 16900 14448 16964 14512
rect 16980 14448 17044 14512
rect 17060 14508 17124 14512
rect 17140 14508 17204 14512
rect 17060 14452 17100 14508
rect 17100 14452 17124 14508
rect 17140 14452 17156 14508
rect 17156 14452 17204 14508
rect 17060 14448 17124 14452
rect 17140 14448 17204 14452
rect 17220 14448 17284 14512
rect 22740 14448 22804 14512
rect 22820 14508 22884 14512
rect 22900 14508 22964 14512
rect 22820 14452 22880 14508
rect 22880 14452 22884 14508
rect 22900 14452 22936 14508
rect 22936 14452 22964 14508
rect 22820 14448 22884 14452
rect 22900 14448 22964 14452
rect 22980 14448 23044 14512
rect 23060 14448 23124 14512
rect 23140 14448 23204 14512
rect 23220 14448 23284 14512
rect 28740 14448 28804 14512
rect 28820 14448 28884 14512
rect 28900 14448 28964 14512
rect 28980 14448 29044 14512
rect 29060 14448 29124 14512
rect 29140 14448 29204 14512
rect 29220 14448 29284 14512
rect 34740 14448 34804 14512
rect 34820 14448 34884 14512
rect 34900 14448 34964 14512
rect 34980 14448 35044 14512
rect 35060 14448 35124 14512
rect 35140 14448 35204 14512
rect 35220 14448 35284 14512
rect 40740 14448 40804 14512
rect 40820 14448 40884 14512
rect 40900 14448 40964 14512
rect 40980 14448 41044 14512
rect 41060 14448 41124 14512
rect 41140 14448 41204 14512
rect 41220 14448 41284 14512
rect 46740 14448 46804 14512
rect 46820 14448 46884 14512
rect 46900 14448 46964 14512
rect 46980 14448 47044 14512
rect 47060 14448 47124 14512
rect 47140 14448 47204 14512
rect 47220 14448 47284 14512
rect 52740 14448 52804 14512
rect 52820 14448 52884 14512
rect 52900 14448 52964 14512
rect 52980 14448 53044 14512
rect 53060 14448 53124 14512
rect 53140 14448 53204 14512
rect 53220 14448 53284 14512
rect 58740 14448 58804 14512
rect 58820 14448 58884 14512
rect 58900 14448 58964 14512
rect 58980 14448 59044 14512
rect 59060 14508 59124 14512
rect 59060 14452 59104 14508
rect 59104 14452 59124 14508
rect 59060 14448 59124 14452
rect 59140 14448 59204 14512
rect 59220 14448 59284 14512
rect 64740 14448 64804 14512
rect 64820 14448 64884 14512
rect 64900 14448 64964 14512
rect 64980 14448 65044 14512
rect 65060 14448 65124 14512
rect 65140 14448 65204 14512
rect 65220 14448 65284 14512
rect 70740 14448 70804 14512
rect 70820 14448 70884 14512
rect 70900 14448 70964 14512
rect 70980 14448 71044 14512
rect 71060 14448 71124 14512
rect 71140 14448 71204 14512
rect 71220 14448 71284 14512
rect 4740 14368 4804 14432
rect 4820 14368 4884 14432
rect 4900 14368 4964 14432
rect 4980 14368 5044 14432
rect 5060 14368 5124 14432
rect 5140 14368 5204 14432
rect 5220 14368 5284 14432
rect 10740 14368 10804 14432
rect 10820 14368 10884 14432
rect 10900 14368 10964 14432
rect 10980 14368 11044 14432
rect 11060 14368 11124 14432
rect 11140 14368 11204 14432
rect 11220 14368 11284 14432
rect 16740 14368 16804 14432
rect 16820 14368 16884 14432
rect 16900 14368 16964 14432
rect 16980 14368 17044 14432
rect 17060 14428 17124 14432
rect 17140 14428 17204 14432
rect 17060 14372 17100 14428
rect 17100 14372 17124 14428
rect 17140 14372 17156 14428
rect 17156 14372 17204 14428
rect 17060 14368 17124 14372
rect 17140 14368 17204 14372
rect 17220 14368 17284 14432
rect 22740 14368 22804 14432
rect 22820 14428 22884 14432
rect 22900 14428 22964 14432
rect 22820 14372 22880 14428
rect 22880 14372 22884 14428
rect 22900 14372 22936 14428
rect 22936 14372 22964 14428
rect 22820 14368 22884 14372
rect 22900 14368 22964 14372
rect 22980 14368 23044 14432
rect 23060 14368 23124 14432
rect 23140 14368 23204 14432
rect 23220 14368 23284 14432
rect 28740 14368 28804 14432
rect 28820 14368 28884 14432
rect 28900 14368 28964 14432
rect 28980 14368 29044 14432
rect 29060 14368 29124 14432
rect 29140 14368 29204 14432
rect 29220 14368 29284 14432
rect 34740 14368 34804 14432
rect 34820 14368 34884 14432
rect 34900 14368 34964 14432
rect 34980 14368 35044 14432
rect 35060 14368 35124 14432
rect 35140 14368 35204 14432
rect 35220 14368 35284 14432
rect 40740 14368 40804 14432
rect 40820 14368 40884 14432
rect 40900 14368 40964 14432
rect 40980 14368 41044 14432
rect 41060 14368 41124 14432
rect 41140 14368 41204 14432
rect 41220 14368 41284 14432
rect 46740 14368 46804 14432
rect 46820 14368 46884 14432
rect 46900 14368 46964 14432
rect 46980 14368 47044 14432
rect 47060 14368 47124 14432
rect 47140 14368 47204 14432
rect 47220 14368 47284 14432
rect 52740 14368 52804 14432
rect 52820 14368 52884 14432
rect 52900 14368 52964 14432
rect 52980 14368 53044 14432
rect 53060 14368 53124 14432
rect 53140 14368 53204 14432
rect 53220 14368 53284 14432
rect 58740 14368 58804 14432
rect 58820 14368 58884 14432
rect 58900 14368 58964 14432
rect 58980 14368 59044 14432
rect 59060 14428 59124 14432
rect 59060 14372 59104 14428
rect 59104 14372 59124 14428
rect 59060 14368 59124 14372
rect 59140 14368 59204 14432
rect 59220 14368 59284 14432
rect 64740 14368 64804 14432
rect 64820 14368 64884 14432
rect 64900 14368 64964 14432
rect 64980 14368 65044 14432
rect 65060 14368 65124 14432
rect 65140 14368 65204 14432
rect 65220 14368 65284 14432
rect 70740 14368 70804 14432
rect 70820 14368 70884 14432
rect 70900 14368 70964 14432
rect 70980 14368 71044 14432
rect 71060 14368 71124 14432
rect 71140 14368 71204 14432
rect 71220 14368 71284 14432
rect 4740 14288 4804 14352
rect 4820 14288 4884 14352
rect 4900 14288 4964 14352
rect 4980 14288 5044 14352
rect 5060 14288 5124 14352
rect 5140 14288 5204 14352
rect 5220 14288 5284 14352
rect 10740 14288 10804 14352
rect 10820 14288 10884 14352
rect 10900 14288 10964 14352
rect 10980 14288 11044 14352
rect 11060 14288 11124 14352
rect 11140 14288 11204 14352
rect 11220 14288 11284 14352
rect 16740 14288 16804 14352
rect 16820 14288 16884 14352
rect 16900 14288 16964 14352
rect 16980 14288 17044 14352
rect 17060 14348 17124 14352
rect 17140 14348 17204 14352
rect 17060 14292 17100 14348
rect 17100 14292 17124 14348
rect 17140 14292 17156 14348
rect 17156 14292 17204 14348
rect 17060 14288 17124 14292
rect 17140 14288 17204 14292
rect 17220 14288 17284 14352
rect 22740 14288 22804 14352
rect 22820 14348 22884 14352
rect 22900 14348 22964 14352
rect 22820 14292 22880 14348
rect 22880 14292 22884 14348
rect 22900 14292 22936 14348
rect 22936 14292 22964 14348
rect 22820 14288 22884 14292
rect 22900 14288 22964 14292
rect 22980 14288 23044 14352
rect 23060 14288 23124 14352
rect 23140 14288 23204 14352
rect 23220 14288 23284 14352
rect 28740 14288 28804 14352
rect 28820 14288 28884 14352
rect 28900 14288 28964 14352
rect 28980 14288 29044 14352
rect 29060 14288 29124 14352
rect 29140 14288 29204 14352
rect 29220 14288 29284 14352
rect 34740 14288 34804 14352
rect 34820 14288 34884 14352
rect 34900 14288 34964 14352
rect 34980 14288 35044 14352
rect 35060 14288 35124 14352
rect 35140 14288 35204 14352
rect 35220 14288 35284 14352
rect 40740 14288 40804 14352
rect 40820 14288 40884 14352
rect 40900 14288 40964 14352
rect 40980 14288 41044 14352
rect 41060 14288 41124 14352
rect 41140 14288 41204 14352
rect 41220 14288 41284 14352
rect 46740 14288 46804 14352
rect 46820 14288 46884 14352
rect 46900 14288 46964 14352
rect 46980 14288 47044 14352
rect 47060 14288 47124 14352
rect 47140 14288 47204 14352
rect 47220 14288 47284 14352
rect 52740 14288 52804 14352
rect 52820 14288 52884 14352
rect 52900 14288 52964 14352
rect 52980 14288 53044 14352
rect 53060 14288 53124 14352
rect 53140 14288 53204 14352
rect 53220 14288 53284 14352
rect 58740 14288 58804 14352
rect 58820 14288 58884 14352
rect 58900 14288 58964 14352
rect 58980 14288 59044 14352
rect 59060 14348 59124 14352
rect 59060 14292 59104 14348
rect 59104 14292 59124 14348
rect 59060 14288 59124 14292
rect 59140 14288 59204 14352
rect 59220 14288 59284 14352
rect 64740 14288 64804 14352
rect 64820 14288 64884 14352
rect 64900 14288 64964 14352
rect 64980 14288 65044 14352
rect 65060 14288 65124 14352
rect 65140 14288 65204 14352
rect 65220 14288 65284 14352
rect 70740 14288 70804 14352
rect 70820 14288 70884 14352
rect 70900 14288 70964 14352
rect 70980 14288 71044 14352
rect 71060 14288 71124 14352
rect 71140 14288 71204 14352
rect 71220 14288 71284 14352
rect 63724 12412 63788 12476
rect 1740 12176 1804 12240
rect 1820 12176 1884 12240
rect 1900 12176 1964 12240
rect 1980 12176 2044 12240
rect 2060 12176 2124 12240
rect 2140 12236 2204 12240
rect 2220 12236 2284 12240
rect 2140 12180 2184 12236
rect 2184 12180 2204 12236
rect 2220 12180 2240 12236
rect 2240 12180 2264 12236
rect 2264 12180 2284 12236
rect 2140 12176 2204 12180
rect 2220 12176 2284 12180
rect 7740 12176 7804 12240
rect 7820 12176 7884 12240
rect 7900 12176 7964 12240
rect 7980 12176 8044 12240
rect 8060 12176 8124 12240
rect 8140 12176 8204 12240
rect 8220 12236 8284 12240
rect 8220 12180 8283 12236
rect 8283 12180 8284 12236
rect 8220 12176 8284 12180
rect 13740 12176 13804 12240
rect 13820 12176 13884 12240
rect 13900 12176 13964 12240
rect 13980 12176 14044 12240
rect 14060 12236 14124 12240
rect 14060 12180 14063 12236
rect 14063 12180 14119 12236
rect 14119 12180 14124 12236
rect 14060 12176 14124 12180
rect 14140 12176 14204 12240
rect 14220 12176 14284 12240
rect 19740 12176 19804 12240
rect 19820 12236 19884 12240
rect 19820 12180 19843 12236
rect 19843 12180 19884 12236
rect 19820 12176 19884 12180
rect 19900 12176 19964 12240
rect 19980 12176 20044 12240
rect 20060 12176 20124 12240
rect 20140 12176 20204 12240
rect 20220 12176 20284 12240
rect 25740 12176 25804 12240
rect 25820 12176 25884 12240
rect 25900 12176 25964 12240
rect 25980 12176 26044 12240
rect 26060 12176 26124 12240
rect 26140 12176 26204 12240
rect 26220 12176 26284 12240
rect 31740 12176 31804 12240
rect 31820 12176 31884 12240
rect 31900 12176 31964 12240
rect 31980 12176 32044 12240
rect 32060 12176 32124 12240
rect 32140 12176 32204 12240
rect 32220 12176 32284 12240
rect 37740 12176 37804 12240
rect 37820 12176 37884 12240
rect 37900 12176 37964 12240
rect 37980 12176 38044 12240
rect 38060 12176 38124 12240
rect 38140 12176 38204 12240
rect 38220 12176 38284 12240
rect 43740 12176 43804 12240
rect 43820 12176 43884 12240
rect 43900 12176 43964 12240
rect 43980 12176 44044 12240
rect 44060 12176 44124 12240
rect 44140 12176 44204 12240
rect 44220 12176 44284 12240
rect 49740 12236 49804 12240
rect 49740 12180 49742 12236
rect 49742 12180 49798 12236
rect 49798 12180 49804 12236
rect 49740 12176 49804 12180
rect 49820 12176 49884 12240
rect 49900 12176 49964 12240
rect 49980 12176 50044 12240
rect 50060 12176 50124 12240
rect 50140 12176 50204 12240
rect 50220 12176 50284 12240
rect 55740 12176 55804 12240
rect 55820 12176 55884 12240
rect 55900 12176 55964 12240
rect 55980 12176 56044 12240
rect 56060 12176 56124 12240
rect 56140 12176 56204 12240
rect 56220 12176 56284 12240
rect 61740 12176 61804 12240
rect 61820 12176 61884 12240
rect 61900 12176 61964 12240
rect 61980 12176 62044 12240
rect 62060 12176 62124 12240
rect 62140 12176 62204 12240
rect 62220 12176 62284 12240
rect 67740 12176 67804 12240
rect 67820 12176 67884 12240
rect 67900 12176 67964 12240
rect 67980 12176 68044 12240
rect 68060 12176 68124 12240
rect 68140 12176 68204 12240
rect 68220 12176 68284 12240
rect 73740 12176 73804 12240
rect 73820 12176 73884 12240
rect 73900 12176 73964 12240
rect 73980 12176 74044 12240
rect 74060 12176 74124 12240
rect 74140 12176 74204 12240
rect 74220 12176 74284 12240
rect 1740 12096 1804 12160
rect 1820 12096 1884 12160
rect 1900 12096 1964 12160
rect 1980 12096 2044 12160
rect 2060 12096 2124 12160
rect 2140 12156 2204 12160
rect 2220 12156 2284 12160
rect 2140 12100 2184 12156
rect 2184 12100 2204 12156
rect 2220 12100 2240 12156
rect 2240 12100 2264 12156
rect 2264 12100 2284 12156
rect 2140 12096 2204 12100
rect 2220 12096 2284 12100
rect 7740 12096 7804 12160
rect 7820 12096 7884 12160
rect 7900 12096 7964 12160
rect 7980 12096 8044 12160
rect 8060 12096 8124 12160
rect 8140 12096 8204 12160
rect 8220 12156 8284 12160
rect 8220 12100 8283 12156
rect 8283 12100 8284 12156
rect 8220 12096 8284 12100
rect 13740 12096 13804 12160
rect 13820 12096 13884 12160
rect 13900 12096 13964 12160
rect 13980 12096 14044 12160
rect 14060 12156 14124 12160
rect 14060 12100 14063 12156
rect 14063 12100 14119 12156
rect 14119 12100 14124 12156
rect 14060 12096 14124 12100
rect 14140 12096 14204 12160
rect 14220 12096 14284 12160
rect 19740 12096 19804 12160
rect 19820 12156 19884 12160
rect 19820 12100 19843 12156
rect 19843 12100 19884 12156
rect 19820 12096 19884 12100
rect 19900 12096 19964 12160
rect 19980 12096 20044 12160
rect 20060 12096 20124 12160
rect 20140 12096 20204 12160
rect 20220 12096 20284 12160
rect 25740 12096 25804 12160
rect 25820 12096 25884 12160
rect 25900 12096 25964 12160
rect 25980 12096 26044 12160
rect 26060 12096 26124 12160
rect 26140 12096 26204 12160
rect 26220 12096 26284 12160
rect 31740 12096 31804 12160
rect 31820 12096 31884 12160
rect 31900 12096 31964 12160
rect 31980 12096 32044 12160
rect 32060 12096 32124 12160
rect 32140 12096 32204 12160
rect 32220 12096 32284 12160
rect 37740 12096 37804 12160
rect 37820 12096 37884 12160
rect 37900 12096 37964 12160
rect 37980 12096 38044 12160
rect 38060 12096 38124 12160
rect 38140 12096 38204 12160
rect 38220 12096 38284 12160
rect 43740 12096 43804 12160
rect 43820 12096 43884 12160
rect 43900 12096 43964 12160
rect 43980 12096 44044 12160
rect 44060 12096 44124 12160
rect 44140 12096 44204 12160
rect 44220 12096 44284 12160
rect 49740 12156 49804 12160
rect 49740 12100 49742 12156
rect 49742 12100 49798 12156
rect 49798 12100 49804 12156
rect 49740 12096 49804 12100
rect 49820 12096 49884 12160
rect 49900 12096 49964 12160
rect 49980 12096 50044 12160
rect 50060 12096 50124 12160
rect 50140 12096 50204 12160
rect 50220 12096 50284 12160
rect 55740 12096 55804 12160
rect 55820 12096 55884 12160
rect 55900 12096 55964 12160
rect 55980 12096 56044 12160
rect 56060 12096 56124 12160
rect 56140 12096 56204 12160
rect 56220 12096 56284 12160
rect 61740 12096 61804 12160
rect 61820 12096 61884 12160
rect 61900 12096 61964 12160
rect 61980 12096 62044 12160
rect 62060 12096 62124 12160
rect 62140 12096 62204 12160
rect 62220 12096 62284 12160
rect 67740 12096 67804 12160
rect 67820 12096 67884 12160
rect 67900 12096 67964 12160
rect 67980 12096 68044 12160
rect 68060 12096 68124 12160
rect 68140 12096 68204 12160
rect 68220 12096 68284 12160
rect 73740 12096 73804 12160
rect 73820 12096 73884 12160
rect 73900 12096 73964 12160
rect 73980 12096 74044 12160
rect 74060 12096 74124 12160
rect 74140 12096 74204 12160
rect 74220 12096 74284 12160
rect 1740 12016 1804 12080
rect 1820 12016 1884 12080
rect 1900 12016 1964 12080
rect 1980 12016 2044 12080
rect 2060 12016 2124 12080
rect 2140 12076 2204 12080
rect 2220 12076 2284 12080
rect 2140 12020 2184 12076
rect 2184 12020 2204 12076
rect 2220 12020 2240 12076
rect 2240 12020 2264 12076
rect 2264 12020 2284 12076
rect 2140 12016 2204 12020
rect 2220 12016 2284 12020
rect 7740 12016 7804 12080
rect 7820 12016 7884 12080
rect 7900 12016 7964 12080
rect 7980 12016 8044 12080
rect 8060 12016 8124 12080
rect 8140 12016 8204 12080
rect 8220 12076 8284 12080
rect 8220 12020 8283 12076
rect 8283 12020 8284 12076
rect 8220 12016 8284 12020
rect 13740 12016 13804 12080
rect 13820 12016 13884 12080
rect 13900 12016 13964 12080
rect 13980 12016 14044 12080
rect 14060 12076 14124 12080
rect 14060 12020 14063 12076
rect 14063 12020 14119 12076
rect 14119 12020 14124 12076
rect 14060 12016 14124 12020
rect 14140 12016 14204 12080
rect 14220 12016 14284 12080
rect 19740 12016 19804 12080
rect 19820 12076 19884 12080
rect 19820 12020 19843 12076
rect 19843 12020 19884 12076
rect 19820 12016 19884 12020
rect 19900 12016 19964 12080
rect 19980 12016 20044 12080
rect 20060 12016 20124 12080
rect 20140 12016 20204 12080
rect 20220 12016 20284 12080
rect 25740 12016 25804 12080
rect 25820 12016 25884 12080
rect 25900 12016 25964 12080
rect 25980 12016 26044 12080
rect 26060 12016 26124 12080
rect 26140 12016 26204 12080
rect 26220 12016 26284 12080
rect 31740 12016 31804 12080
rect 31820 12016 31884 12080
rect 31900 12016 31964 12080
rect 31980 12016 32044 12080
rect 32060 12016 32124 12080
rect 32140 12016 32204 12080
rect 32220 12016 32284 12080
rect 37740 12016 37804 12080
rect 37820 12016 37884 12080
rect 37900 12016 37964 12080
rect 37980 12016 38044 12080
rect 38060 12016 38124 12080
rect 38140 12016 38204 12080
rect 38220 12016 38284 12080
rect 43740 12016 43804 12080
rect 43820 12016 43884 12080
rect 43900 12016 43964 12080
rect 43980 12016 44044 12080
rect 44060 12016 44124 12080
rect 44140 12016 44204 12080
rect 44220 12016 44284 12080
rect 49740 12076 49804 12080
rect 49740 12020 49742 12076
rect 49742 12020 49798 12076
rect 49798 12020 49804 12076
rect 49740 12016 49804 12020
rect 49820 12016 49884 12080
rect 49900 12016 49964 12080
rect 49980 12016 50044 12080
rect 50060 12016 50124 12080
rect 50140 12016 50204 12080
rect 50220 12016 50284 12080
rect 55740 12016 55804 12080
rect 55820 12016 55884 12080
rect 55900 12016 55964 12080
rect 55980 12016 56044 12080
rect 56060 12016 56124 12080
rect 56140 12016 56204 12080
rect 56220 12016 56284 12080
rect 61740 12016 61804 12080
rect 61820 12016 61884 12080
rect 61900 12016 61964 12080
rect 61980 12016 62044 12080
rect 62060 12016 62124 12080
rect 62140 12016 62204 12080
rect 62220 12016 62284 12080
rect 67740 12016 67804 12080
rect 67820 12016 67884 12080
rect 67900 12016 67964 12080
rect 67980 12016 68044 12080
rect 68060 12016 68124 12080
rect 68140 12016 68204 12080
rect 68220 12016 68284 12080
rect 73740 12016 73804 12080
rect 73820 12016 73884 12080
rect 73900 12016 73964 12080
rect 73980 12016 74044 12080
rect 74060 12016 74124 12080
rect 74140 12016 74204 12080
rect 74220 12016 74284 12080
rect 1740 11936 1804 12000
rect 1820 11936 1884 12000
rect 1900 11936 1964 12000
rect 1980 11936 2044 12000
rect 2060 11936 2124 12000
rect 2140 11996 2204 12000
rect 2220 11996 2284 12000
rect 2140 11940 2184 11996
rect 2184 11940 2204 11996
rect 2220 11940 2240 11996
rect 2240 11940 2264 11996
rect 2264 11940 2284 11996
rect 2140 11936 2204 11940
rect 2220 11936 2284 11940
rect 7740 11936 7804 12000
rect 7820 11936 7884 12000
rect 7900 11936 7964 12000
rect 7980 11936 8044 12000
rect 8060 11936 8124 12000
rect 8140 11936 8204 12000
rect 8220 11996 8284 12000
rect 8220 11940 8283 11996
rect 8283 11940 8284 11996
rect 8220 11936 8284 11940
rect 13740 11936 13804 12000
rect 13820 11936 13884 12000
rect 13900 11936 13964 12000
rect 13980 11936 14044 12000
rect 14060 11996 14124 12000
rect 14060 11940 14063 11996
rect 14063 11940 14119 11996
rect 14119 11940 14124 11996
rect 14060 11936 14124 11940
rect 14140 11936 14204 12000
rect 14220 11936 14284 12000
rect 19740 11936 19804 12000
rect 19820 11996 19884 12000
rect 19820 11940 19843 11996
rect 19843 11940 19884 11996
rect 19820 11936 19884 11940
rect 19900 11936 19964 12000
rect 19980 11936 20044 12000
rect 20060 11936 20124 12000
rect 20140 11936 20204 12000
rect 20220 11936 20284 12000
rect 25740 11936 25804 12000
rect 25820 11936 25884 12000
rect 25900 11936 25964 12000
rect 25980 11936 26044 12000
rect 26060 11936 26124 12000
rect 26140 11936 26204 12000
rect 26220 11936 26284 12000
rect 31740 11936 31804 12000
rect 31820 11936 31884 12000
rect 31900 11936 31964 12000
rect 31980 11936 32044 12000
rect 32060 11936 32124 12000
rect 32140 11936 32204 12000
rect 32220 11936 32284 12000
rect 37740 11936 37804 12000
rect 37820 11936 37884 12000
rect 37900 11936 37964 12000
rect 37980 11936 38044 12000
rect 38060 11936 38124 12000
rect 38140 11936 38204 12000
rect 38220 11936 38284 12000
rect 43740 11936 43804 12000
rect 43820 11936 43884 12000
rect 43900 11936 43964 12000
rect 43980 11936 44044 12000
rect 44060 11936 44124 12000
rect 44140 11936 44204 12000
rect 44220 11936 44284 12000
rect 49740 11996 49804 12000
rect 49740 11940 49742 11996
rect 49742 11940 49798 11996
rect 49798 11940 49804 11996
rect 49740 11936 49804 11940
rect 49820 11936 49884 12000
rect 49900 11936 49964 12000
rect 49980 11936 50044 12000
rect 50060 11936 50124 12000
rect 50140 11936 50204 12000
rect 50220 11936 50284 12000
rect 55740 11936 55804 12000
rect 55820 11936 55884 12000
rect 55900 11936 55964 12000
rect 55980 11936 56044 12000
rect 56060 11936 56124 12000
rect 56140 11936 56204 12000
rect 56220 11936 56284 12000
rect 61740 11936 61804 12000
rect 61820 11936 61884 12000
rect 61900 11936 61964 12000
rect 61980 11936 62044 12000
rect 62060 11936 62124 12000
rect 62140 11936 62204 12000
rect 62220 11936 62284 12000
rect 67740 11936 67804 12000
rect 67820 11936 67884 12000
rect 67900 11936 67964 12000
rect 67980 11936 68044 12000
rect 68060 11936 68124 12000
rect 68140 11936 68204 12000
rect 68220 11936 68284 12000
rect 73740 11936 73804 12000
rect 73820 11936 73884 12000
rect 73900 11936 73964 12000
rect 73980 11936 74044 12000
rect 74060 11936 74124 12000
rect 74140 11936 74204 12000
rect 74220 11936 74284 12000
rect 63724 11792 63788 11796
rect 63724 11736 63738 11792
rect 63738 11736 63788 11792
rect 63724 11732 63788 11736
rect 65564 11596 65628 11660
rect 66116 11596 66180 11660
rect 65564 11460 65628 11524
rect 63908 7652 63972 7716
rect 65564 7652 65628 7716
rect 65748 7516 65812 7580
rect 62988 6896 63052 6900
rect 62988 6840 63002 6896
rect 63002 6840 63052 6896
rect 62988 6836 63052 6840
rect 66668 6836 66732 6900
rect 64460 6700 64524 6764
rect 65932 6156 65996 6220
rect 39988 5748 40052 5812
rect 68508 5612 68572 5676
rect 64092 5340 64156 5404
rect 66484 5204 66548 5268
rect 64276 4932 64340 4996
rect 63172 4796 63236 4860
rect 4740 4528 4804 4592
rect 4820 4528 4884 4592
rect 4900 4528 4964 4592
rect 4980 4528 5044 4592
rect 5060 4528 5124 4592
rect 5140 4528 5204 4592
rect 5220 4528 5284 4592
rect 10740 4528 10804 4592
rect 10820 4528 10884 4592
rect 10900 4528 10964 4592
rect 10980 4528 11044 4592
rect 11060 4528 11124 4592
rect 11140 4528 11204 4592
rect 11220 4528 11284 4592
rect 16740 4528 16804 4592
rect 16820 4528 16884 4592
rect 16900 4528 16964 4592
rect 16980 4528 17044 4592
rect 17060 4528 17124 4592
rect 17140 4528 17204 4592
rect 17220 4528 17284 4592
rect 22740 4528 22804 4592
rect 22820 4528 22884 4592
rect 22900 4528 22964 4592
rect 22980 4528 23044 4592
rect 23060 4528 23124 4592
rect 23140 4528 23204 4592
rect 23220 4528 23284 4592
rect 28740 4528 28804 4592
rect 28820 4528 28884 4592
rect 28900 4528 28964 4592
rect 28980 4528 29044 4592
rect 29060 4528 29124 4592
rect 29140 4528 29204 4592
rect 29220 4528 29284 4592
rect 34740 4528 34804 4592
rect 34820 4528 34884 4592
rect 34900 4528 34964 4592
rect 34980 4528 35044 4592
rect 35060 4528 35124 4592
rect 35140 4528 35204 4592
rect 35220 4528 35284 4592
rect 40740 4528 40804 4592
rect 40820 4528 40884 4592
rect 40900 4528 40964 4592
rect 40980 4528 41044 4592
rect 41060 4528 41124 4592
rect 41140 4528 41204 4592
rect 41220 4528 41284 4592
rect 46740 4528 46804 4592
rect 46820 4528 46884 4592
rect 46900 4528 46964 4592
rect 46980 4528 47044 4592
rect 47060 4528 47124 4592
rect 47140 4528 47204 4592
rect 47220 4528 47284 4592
rect 52740 4528 52804 4592
rect 52820 4528 52884 4592
rect 52900 4528 52964 4592
rect 52980 4528 53044 4592
rect 53060 4528 53124 4592
rect 53140 4528 53204 4592
rect 53220 4528 53284 4592
rect 58740 4528 58804 4592
rect 58820 4528 58884 4592
rect 58900 4528 58964 4592
rect 58980 4528 59044 4592
rect 59060 4528 59124 4592
rect 59140 4528 59204 4592
rect 59220 4528 59284 4592
rect 64740 4528 64804 4592
rect 64820 4528 64884 4592
rect 64900 4528 64964 4592
rect 64980 4528 65044 4592
rect 65060 4528 65124 4592
rect 65140 4528 65204 4592
rect 65220 4528 65284 4592
rect 70740 4528 70804 4592
rect 70820 4528 70884 4592
rect 70900 4528 70964 4592
rect 70980 4528 71044 4592
rect 71060 4528 71124 4592
rect 71140 4528 71204 4592
rect 71220 4528 71284 4592
rect 4740 4448 4804 4512
rect 4820 4448 4884 4512
rect 4900 4448 4964 4512
rect 4980 4448 5044 4512
rect 5060 4448 5124 4512
rect 5140 4448 5204 4512
rect 5220 4448 5284 4512
rect 10740 4448 10804 4512
rect 10820 4448 10884 4512
rect 10900 4448 10964 4512
rect 10980 4448 11044 4512
rect 11060 4448 11124 4512
rect 11140 4448 11204 4512
rect 11220 4448 11284 4512
rect 16740 4448 16804 4512
rect 16820 4448 16884 4512
rect 16900 4448 16964 4512
rect 16980 4448 17044 4512
rect 17060 4448 17124 4512
rect 17140 4448 17204 4512
rect 17220 4448 17284 4512
rect 22740 4448 22804 4512
rect 22820 4448 22884 4512
rect 22900 4448 22964 4512
rect 22980 4448 23044 4512
rect 23060 4448 23124 4512
rect 23140 4448 23204 4512
rect 23220 4448 23284 4512
rect 28740 4448 28804 4512
rect 28820 4448 28884 4512
rect 28900 4448 28964 4512
rect 28980 4448 29044 4512
rect 29060 4448 29124 4512
rect 29140 4448 29204 4512
rect 29220 4448 29284 4512
rect 34740 4448 34804 4512
rect 34820 4448 34884 4512
rect 34900 4448 34964 4512
rect 34980 4448 35044 4512
rect 35060 4448 35124 4512
rect 35140 4448 35204 4512
rect 35220 4448 35284 4512
rect 40740 4448 40804 4512
rect 40820 4448 40884 4512
rect 40900 4448 40964 4512
rect 40980 4448 41044 4512
rect 41060 4448 41124 4512
rect 41140 4448 41204 4512
rect 41220 4448 41284 4512
rect 46740 4448 46804 4512
rect 46820 4448 46884 4512
rect 46900 4448 46964 4512
rect 46980 4448 47044 4512
rect 47060 4448 47124 4512
rect 47140 4448 47204 4512
rect 47220 4448 47284 4512
rect 52740 4448 52804 4512
rect 52820 4448 52884 4512
rect 52900 4448 52964 4512
rect 52980 4448 53044 4512
rect 53060 4448 53124 4512
rect 53140 4448 53204 4512
rect 53220 4448 53284 4512
rect 58740 4448 58804 4512
rect 58820 4448 58884 4512
rect 58900 4448 58964 4512
rect 58980 4448 59044 4512
rect 59060 4448 59124 4512
rect 59140 4448 59204 4512
rect 59220 4448 59284 4512
rect 64740 4448 64804 4512
rect 64820 4448 64884 4512
rect 64900 4448 64964 4512
rect 64980 4448 65044 4512
rect 65060 4448 65124 4512
rect 65140 4448 65204 4512
rect 65220 4448 65284 4512
rect 70740 4448 70804 4512
rect 70820 4448 70884 4512
rect 70900 4448 70964 4512
rect 70980 4448 71044 4512
rect 71060 4448 71124 4512
rect 71140 4448 71204 4512
rect 71220 4448 71284 4512
rect 4740 4368 4804 4432
rect 4820 4368 4884 4432
rect 4900 4368 4964 4432
rect 4980 4368 5044 4432
rect 5060 4368 5124 4432
rect 5140 4368 5204 4432
rect 5220 4368 5284 4432
rect 10740 4368 10804 4432
rect 10820 4368 10884 4432
rect 10900 4368 10964 4432
rect 10980 4368 11044 4432
rect 11060 4368 11124 4432
rect 11140 4368 11204 4432
rect 11220 4368 11284 4432
rect 16740 4368 16804 4432
rect 16820 4368 16884 4432
rect 16900 4368 16964 4432
rect 16980 4368 17044 4432
rect 17060 4368 17124 4432
rect 17140 4368 17204 4432
rect 17220 4368 17284 4432
rect 22740 4368 22804 4432
rect 22820 4368 22884 4432
rect 22900 4368 22964 4432
rect 22980 4368 23044 4432
rect 23060 4368 23124 4432
rect 23140 4368 23204 4432
rect 23220 4368 23284 4432
rect 28740 4368 28804 4432
rect 28820 4368 28884 4432
rect 28900 4368 28964 4432
rect 28980 4368 29044 4432
rect 29060 4368 29124 4432
rect 29140 4368 29204 4432
rect 29220 4368 29284 4432
rect 34740 4368 34804 4432
rect 34820 4368 34884 4432
rect 34900 4368 34964 4432
rect 34980 4368 35044 4432
rect 35060 4368 35124 4432
rect 35140 4368 35204 4432
rect 35220 4368 35284 4432
rect 40740 4368 40804 4432
rect 40820 4368 40884 4432
rect 40900 4368 40964 4432
rect 40980 4368 41044 4432
rect 41060 4368 41124 4432
rect 41140 4368 41204 4432
rect 41220 4368 41284 4432
rect 46740 4368 46804 4432
rect 46820 4368 46884 4432
rect 46900 4368 46964 4432
rect 46980 4368 47044 4432
rect 47060 4368 47124 4432
rect 47140 4368 47204 4432
rect 47220 4368 47284 4432
rect 52740 4368 52804 4432
rect 52820 4368 52884 4432
rect 52900 4368 52964 4432
rect 52980 4368 53044 4432
rect 53060 4368 53124 4432
rect 53140 4368 53204 4432
rect 53220 4368 53284 4432
rect 58740 4368 58804 4432
rect 58820 4368 58884 4432
rect 58900 4368 58964 4432
rect 58980 4368 59044 4432
rect 59060 4368 59124 4432
rect 59140 4368 59204 4432
rect 59220 4368 59284 4432
rect 64740 4368 64804 4432
rect 64820 4368 64884 4432
rect 64900 4368 64964 4432
rect 64980 4368 65044 4432
rect 65060 4368 65124 4432
rect 65140 4368 65204 4432
rect 65220 4368 65284 4432
rect 70740 4368 70804 4432
rect 70820 4368 70884 4432
rect 70900 4368 70964 4432
rect 70980 4368 71044 4432
rect 71060 4368 71124 4432
rect 71140 4368 71204 4432
rect 71220 4368 71284 4432
rect 4740 4288 4804 4352
rect 4820 4288 4884 4352
rect 4900 4288 4964 4352
rect 4980 4288 5044 4352
rect 5060 4288 5124 4352
rect 5140 4288 5204 4352
rect 5220 4288 5284 4352
rect 10740 4288 10804 4352
rect 10820 4288 10884 4352
rect 10900 4288 10964 4352
rect 10980 4288 11044 4352
rect 11060 4288 11124 4352
rect 11140 4288 11204 4352
rect 11220 4288 11284 4352
rect 16740 4288 16804 4352
rect 16820 4288 16884 4352
rect 16900 4288 16964 4352
rect 16980 4288 17044 4352
rect 17060 4288 17124 4352
rect 17140 4288 17204 4352
rect 17220 4288 17284 4352
rect 22740 4288 22804 4352
rect 22820 4288 22884 4352
rect 22900 4288 22964 4352
rect 22980 4288 23044 4352
rect 23060 4288 23124 4352
rect 23140 4288 23204 4352
rect 23220 4288 23284 4352
rect 28740 4288 28804 4352
rect 28820 4288 28884 4352
rect 28900 4288 28964 4352
rect 28980 4288 29044 4352
rect 29060 4288 29124 4352
rect 29140 4288 29204 4352
rect 29220 4288 29284 4352
rect 34740 4288 34804 4352
rect 34820 4288 34884 4352
rect 34900 4288 34964 4352
rect 34980 4288 35044 4352
rect 35060 4288 35124 4352
rect 35140 4288 35204 4352
rect 35220 4288 35284 4352
rect 40740 4288 40804 4352
rect 40820 4288 40884 4352
rect 40900 4288 40964 4352
rect 40980 4288 41044 4352
rect 41060 4288 41124 4352
rect 41140 4288 41204 4352
rect 41220 4288 41284 4352
rect 46740 4288 46804 4352
rect 46820 4288 46884 4352
rect 46900 4288 46964 4352
rect 46980 4288 47044 4352
rect 47060 4288 47124 4352
rect 47140 4288 47204 4352
rect 47220 4288 47284 4352
rect 52740 4288 52804 4352
rect 52820 4288 52884 4352
rect 52900 4288 52964 4352
rect 52980 4288 53044 4352
rect 53060 4288 53124 4352
rect 53140 4288 53204 4352
rect 53220 4288 53284 4352
rect 58740 4288 58804 4352
rect 58820 4288 58884 4352
rect 58900 4288 58964 4352
rect 58980 4288 59044 4352
rect 59060 4288 59124 4352
rect 59140 4288 59204 4352
rect 59220 4288 59284 4352
rect 64740 4288 64804 4352
rect 64820 4288 64884 4352
rect 64900 4288 64964 4352
rect 64980 4288 65044 4352
rect 65060 4288 65124 4352
rect 65140 4288 65204 4352
rect 65220 4288 65284 4352
rect 70740 4288 70804 4352
rect 70820 4288 70884 4352
rect 70900 4288 70964 4352
rect 70980 4288 71044 4352
rect 71060 4288 71124 4352
rect 71140 4288 71204 4352
rect 71220 4288 71284 4352
rect 66116 3980 66180 4044
rect 39988 3300 40052 3364
rect 66300 3300 66364 3364
rect 1740 2176 1804 2240
rect 1820 2236 1884 2240
rect 1900 2236 1964 2240
rect 1980 2236 2044 2240
rect 2060 2236 2124 2240
rect 2140 2236 2204 2240
rect 1820 2180 1864 2236
rect 1864 2180 1884 2236
rect 1900 2180 1920 2236
rect 1920 2180 1944 2236
rect 1944 2180 1964 2236
rect 1980 2180 2000 2236
rect 2000 2180 2024 2236
rect 2024 2180 2044 2236
rect 2060 2180 2080 2236
rect 2080 2180 2104 2236
rect 2104 2180 2124 2236
rect 2140 2180 2160 2236
rect 2160 2180 2204 2236
rect 1820 2176 1884 2180
rect 1900 2176 1964 2180
rect 1980 2176 2044 2180
rect 2060 2176 2124 2180
rect 2140 2176 2204 2180
rect 2220 2176 2284 2240
rect 7740 2176 7804 2240
rect 7820 2176 7884 2240
rect 7900 2176 7964 2240
rect 7980 2176 8044 2240
rect 8060 2176 8124 2240
rect 8140 2176 8204 2240
rect 8220 2176 8284 2240
rect 13740 2176 13804 2240
rect 13820 2176 13884 2240
rect 13900 2176 13964 2240
rect 13980 2176 14044 2240
rect 14060 2176 14124 2240
rect 14140 2176 14204 2240
rect 14220 2176 14284 2240
rect 19740 2176 19804 2240
rect 19820 2176 19884 2240
rect 19900 2176 19964 2240
rect 19980 2176 20044 2240
rect 20060 2176 20124 2240
rect 20140 2176 20204 2240
rect 20220 2176 20284 2240
rect 25740 2176 25804 2240
rect 25820 2176 25884 2240
rect 25900 2176 25964 2240
rect 25980 2176 26044 2240
rect 26060 2176 26124 2240
rect 26140 2176 26204 2240
rect 26220 2176 26284 2240
rect 31740 2176 31804 2240
rect 31820 2236 31884 2240
rect 31900 2236 31964 2240
rect 31980 2236 32044 2240
rect 32060 2236 32124 2240
rect 32140 2236 32204 2240
rect 31820 2180 31864 2236
rect 31864 2180 31884 2236
rect 31900 2180 31920 2236
rect 31920 2180 31944 2236
rect 31944 2180 31964 2236
rect 31980 2180 32000 2236
rect 32000 2180 32024 2236
rect 32024 2180 32044 2236
rect 32060 2180 32080 2236
rect 32080 2180 32104 2236
rect 32104 2180 32124 2236
rect 32140 2180 32160 2236
rect 32160 2180 32204 2236
rect 31820 2176 31884 2180
rect 31900 2176 31964 2180
rect 31980 2176 32044 2180
rect 32060 2176 32124 2180
rect 32140 2176 32204 2180
rect 32220 2176 32284 2240
rect 37740 2176 37804 2240
rect 37820 2176 37884 2240
rect 37900 2176 37964 2240
rect 37980 2176 38044 2240
rect 38060 2176 38124 2240
rect 38140 2176 38204 2240
rect 38220 2176 38284 2240
rect 43740 2176 43804 2240
rect 43820 2176 43884 2240
rect 43900 2176 43964 2240
rect 43980 2176 44044 2240
rect 44060 2176 44124 2240
rect 44140 2176 44204 2240
rect 44220 2176 44284 2240
rect 49740 2176 49804 2240
rect 49820 2176 49884 2240
rect 49900 2176 49964 2240
rect 49980 2176 50044 2240
rect 50060 2176 50124 2240
rect 50140 2176 50204 2240
rect 50220 2176 50284 2240
rect 55740 2176 55804 2240
rect 55820 2176 55884 2240
rect 55900 2176 55964 2240
rect 55980 2176 56044 2240
rect 56060 2176 56124 2240
rect 56140 2176 56204 2240
rect 56220 2176 56284 2240
rect 61740 2176 61804 2240
rect 61820 2236 61884 2240
rect 61900 2236 61964 2240
rect 61980 2236 62044 2240
rect 62060 2236 62124 2240
rect 62140 2236 62204 2240
rect 61820 2180 61864 2236
rect 61864 2180 61884 2236
rect 61900 2180 61920 2236
rect 61920 2180 61944 2236
rect 61944 2180 61964 2236
rect 61980 2180 62000 2236
rect 62000 2180 62024 2236
rect 62024 2180 62044 2236
rect 62060 2180 62080 2236
rect 62080 2180 62104 2236
rect 62104 2180 62124 2236
rect 62140 2180 62160 2236
rect 62160 2180 62204 2236
rect 61820 2176 61884 2180
rect 61900 2176 61964 2180
rect 61980 2176 62044 2180
rect 62060 2176 62124 2180
rect 62140 2176 62204 2180
rect 62220 2176 62284 2240
rect 67740 2176 67804 2240
rect 67820 2176 67884 2240
rect 67900 2176 67964 2240
rect 67980 2176 68044 2240
rect 68060 2176 68124 2240
rect 68140 2176 68204 2240
rect 68220 2176 68284 2240
rect 73740 2176 73804 2240
rect 73820 2176 73884 2240
rect 73900 2176 73964 2240
rect 73980 2176 74044 2240
rect 74060 2176 74124 2240
rect 74140 2176 74204 2240
rect 74220 2176 74284 2240
rect 1740 2096 1804 2160
rect 1820 2156 1884 2160
rect 1900 2156 1964 2160
rect 1980 2156 2044 2160
rect 2060 2156 2124 2160
rect 2140 2156 2204 2160
rect 1820 2100 1864 2156
rect 1864 2100 1884 2156
rect 1900 2100 1920 2156
rect 1920 2100 1944 2156
rect 1944 2100 1964 2156
rect 1980 2100 2000 2156
rect 2000 2100 2024 2156
rect 2024 2100 2044 2156
rect 2060 2100 2080 2156
rect 2080 2100 2104 2156
rect 2104 2100 2124 2156
rect 2140 2100 2160 2156
rect 2160 2100 2204 2156
rect 1820 2096 1884 2100
rect 1900 2096 1964 2100
rect 1980 2096 2044 2100
rect 2060 2096 2124 2100
rect 2140 2096 2204 2100
rect 2220 2096 2284 2160
rect 7740 2096 7804 2160
rect 7820 2096 7884 2160
rect 7900 2096 7964 2160
rect 7980 2096 8044 2160
rect 8060 2096 8124 2160
rect 8140 2096 8204 2160
rect 8220 2096 8284 2160
rect 13740 2096 13804 2160
rect 13820 2096 13884 2160
rect 13900 2096 13964 2160
rect 13980 2096 14044 2160
rect 14060 2096 14124 2160
rect 14140 2096 14204 2160
rect 14220 2096 14284 2160
rect 19740 2096 19804 2160
rect 19820 2096 19884 2160
rect 19900 2096 19964 2160
rect 19980 2096 20044 2160
rect 20060 2096 20124 2160
rect 20140 2096 20204 2160
rect 20220 2096 20284 2160
rect 25740 2096 25804 2160
rect 25820 2096 25884 2160
rect 25900 2096 25964 2160
rect 25980 2096 26044 2160
rect 26060 2096 26124 2160
rect 26140 2096 26204 2160
rect 26220 2096 26284 2160
rect 31740 2096 31804 2160
rect 31820 2156 31884 2160
rect 31900 2156 31964 2160
rect 31980 2156 32044 2160
rect 32060 2156 32124 2160
rect 32140 2156 32204 2160
rect 31820 2100 31864 2156
rect 31864 2100 31884 2156
rect 31900 2100 31920 2156
rect 31920 2100 31944 2156
rect 31944 2100 31964 2156
rect 31980 2100 32000 2156
rect 32000 2100 32024 2156
rect 32024 2100 32044 2156
rect 32060 2100 32080 2156
rect 32080 2100 32104 2156
rect 32104 2100 32124 2156
rect 32140 2100 32160 2156
rect 32160 2100 32204 2156
rect 31820 2096 31884 2100
rect 31900 2096 31964 2100
rect 31980 2096 32044 2100
rect 32060 2096 32124 2100
rect 32140 2096 32204 2100
rect 32220 2096 32284 2160
rect 37740 2096 37804 2160
rect 37820 2096 37884 2160
rect 37900 2096 37964 2160
rect 37980 2096 38044 2160
rect 38060 2096 38124 2160
rect 38140 2096 38204 2160
rect 38220 2096 38284 2160
rect 43740 2096 43804 2160
rect 43820 2096 43884 2160
rect 43900 2096 43964 2160
rect 43980 2096 44044 2160
rect 44060 2096 44124 2160
rect 44140 2096 44204 2160
rect 44220 2096 44284 2160
rect 49740 2096 49804 2160
rect 49820 2096 49884 2160
rect 49900 2096 49964 2160
rect 49980 2096 50044 2160
rect 50060 2096 50124 2160
rect 50140 2096 50204 2160
rect 50220 2096 50284 2160
rect 55740 2096 55804 2160
rect 55820 2096 55884 2160
rect 55900 2096 55964 2160
rect 55980 2096 56044 2160
rect 56060 2096 56124 2160
rect 56140 2096 56204 2160
rect 56220 2096 56284 2160
rect 61740 2096 61804 2160
rect 61820 2156 61884 2160
rect 61900 2156 61964 2160
rect 61980 2156 62044 2160
rect 62060 2156 62124 2160
rect 62140 2156 62204 2160
rect 61820 2100 61864 2156
rect 61864 2100 61884 2156
rect 61900 2100 61920 2156
rect 61920 2100 61944 2156
rect 61944 2100 61964 2156
rect 61980 2100 62000 2156
rect 62000 2100 62024 2156
rect 62024 2100 62044 2156
rect 62060 2100 62080 2156
rect 62080 2100 62104 2156
rect 62104 2100 62124 2156
rect 62140 2100 62160 2156
rect 62160 2100 62204 2156
rect 61820 2096 61884 2100
rect 61900 2096 61964 2100
rect 61980 2096 62044 2100
rect 62060 2096 62124 2100
rect 62140 2096 62204 2100
rect 62220 2096 62284 2160
rect 67740 2096 67804 2160
rect 67820 2096 67884 2160
rect 67900 2096 67964 2160
rect 67980 2096 68044 2160
rect 68060 2096 68124 2160
rect 68140 2096 68204 2160
rect 68220 2096 68284 2160
rect 73740 2096 73804 2160
rect 73820 2096 73884 2160
rect 73900 2096 73964 2160
rect 73980 2096 74044 2160
rect 74060 2096 74124 2160
rect 74140 2096 74204 2160
rect 74220 2096 74284 2160
rect 1740 2016 1804 2080
rect 1820 2076 1884 2080
rect 1900 2076 1964 2080
rect 1980 2076 2044 2080
rect 2060 2076 2124 2080
rect 2140 2076 2204 2080
rect 1820 2020 1864 2076
rect 1864 2020 1884 2076
rect 1900 2020 1920 2076
rect 1920 2020 1944 2076
rect 1944 2020 1964 2076
rect 1980 2020 2000 2076
rect 2000 2020 2024 2076
rect 2024 2020 2044 2076
rect 2060 2020 2080 2076
rect 2080 2020 2104 2076
rect 2104 2020 2124 2076
rect 2140 2020 2160 2076
rect 2160 2020 2204 2076
rect 1820 2016 1884 2020
rect 1900 2016 1964 2020
rect 1980 2016 2044 2020
rect 2060 2016 2124 2020
rect 2140 2016 2204 2020
rect 2220 2016 2284 2080
rect 7740 2016 7804 2080
rect 7820 2016 7884 2080
rect 7900 2016 7964 2080
rect 7980 2016 8044 2080
rect 8060 2016 8124 2080
rect 8140 2016 8204 2080
rect 8220 2016 8284 2080
rect 13740 2016 13804 2080
rect 13820 2016 13884 2080
rect 13900 2016 13964 2080
rect 13980 2016 14044 2080
rect 14060 2016 14124 2080
rect 14140 2016 14204 2080
rect 14220 2016 14284 2080
rect 19740 2016 19804 2080
rect 19820 2016 19884 2080
rect 19900 2016 19964 2080
rect 19980 2016 20044 2080
rect 20060 2016 20124 2080
rect 20140 2016 20204 2080
rect 20220 2016 20284 2080
rect 25740 2016 25804 2080
rect 25820 2016 25884 2080
rect 25900 2016 25964 2080
rect 25980 2016 26044 2080
rect 26060 2016 26124 2080
rect 26140 2016 26204 2080
rect 26220 2016 26284 2080
rect 31740 2016 31804 2080
rect 31820 2076 31884 2080
rect 31900 2076 31964 2080
rect 31980 2076 32044 2080
rect 32060 2076 32124 2080
rect 32140 2076 32204 2080
rect 31820 2020 31864 2076
rect 31864 2020 31884 2076
rect 31900 2020 31920 2076
rect 31920 2020 31944 2076
rect 31944 2020 31964 2076
rect 31980 2020 32000 2076
rect 32000 2020 32024 2076
rect 32024 2020 32044 2076
rect 32060 2020 32080 2076
rect 32080 2020 32104 2076
rect 32104 2020 32124 2076
rect 32140 2020 32160 2076
rect 32160 2020 32204 2076
rect 31820 2016 31884 2020
rect 31900 2016 31964 2020
rect 31980 2016 32044 2020
rect 32060 2016 32124 2020
rect 32140 2016 32204 2020
rect 32220 2016 32284 2080
rect 37740 2016 37804 2080
rect 37820 2016 37884 2080
rect 37900 2016 37964 2080
rect 37980 2016 38044 2080
rect 38060 2016 38124 2080
rect 38140 2016 38204 2080
rect 38220 2016 38284 2080
rect 43740 2016 43804 2080
rect 43820 2016 43884 2080
rect 43900 2016 43964 2080
rect 43980 2016 44044 2080
rect 44060 2016 44124 2080
rect 44140 2016 44204 2080
rect 44220 2016 44284 2080
rect 49740 2016 49804 2080
rect 49820 2016 49884 2080
rect 49900 2016 49964 2080
rect 49980 2016 50044 2080
rect 50060 2016 50124 2080
rect 50140 2016 50204 2080
rect 50220 2016 50284 2080
rect 55740 2016 55804 2080
rect 55820 2016 55884 2080
rect 55900 2016 55964 2080
rect 55980 2016 56044 2080
rect 56060 2016 56124 2080
rect 56140 2016 56204 2080
rect 56220 2016 56284 2080
rect 61740 2016 61804 2080
rect 61820 2076 61884 2080
rect 61900 2076 61964 2080
rect 61980 2076 62044 2080
rect 62060 2076 62124 2080
rect 62140 2076 62204 2080
rect 61820 2020 61864 2076
rect 61864 2020 61884 2076
rect 61900 2020 61920 2076
rect 61920 2020 61944 2076
rect 61944 2020 61964 2076
rect 61980 2020 62000 2076
rect 62000 2020 62024 2076
rect 62024 2020 62044 2076
rect 62060 2020 62080 2076
rect 62080 2020 62104 2076
rect 62104 2020 62124 2076
rect 62140 2020 62160 2076
rect 62160 2020 62204 2076
rect 61820 2016 61884 2020
rect 61900 2016 61964 2020
rect 61980 2016 62044 2020
rect 62060 2016 62124 2020
rect 62140 2016 62204 2020
rect 62220 2016 62284 2080
rect 67740 2016 67804 2080
rect 67820 2016 67884 2080
rect 67900 2016 67964 2080
rect 67980 2016 68044 2080
rect 68060 2016 68124 2080
rect 68140 2016 68204 2080
rect 68220 2016 68284 2080
rect 73740 2016 73804 2080
rect 73820 2016 73884 2080
rect 73900 2016 73964 2080
rect 73980 2016 74044 2080
rect 74060 2016 74124 2080
rect 74140 2016 74204 2080
rect 74220 2016 74284 2080
rect 1740 1936 1804 2000
rect 1820 1996 1884 2000
rect 1900 1996 1964 2000
rect 1980 1996 2044 2000
rect 2060 1996 2124 2000
rect 2140 1996 2204 2000
rect 1820 1940 1864 1996
rect 1864 1940 1884 1996
rect 1900 1940 1920 1996
rect 1920 1940 1944 1996
rect 1944 1940 1964 1996
rect 1980 1940 2000 1996
rect 2000 1940 2024 1996
rect 2024 1940 2044 1996
rect 2060 1940 2080 1996
rect 2080 1940 2104 1996
rect 2104 1940 2124 1996
rect 2140 1940 2160 1996
rect 2160 1940 2204 1996
rect 1820 1936 1884 1940
rect 1900 1936 1964 1940
rect 1980 1936 2044 1940
rect 2060 1936 2124 1940
rect 2140 1936 2204 1940
rect 2220 1936 2284 2000
rect 7740 1936 7804 2000
rect 7820 1936 7884 2000
rect 7900 1936 7964 2000
rect 7980 1936 8044 2000
rect 8060 1936 8124 2000
rect 8140 1936 8204 2000
rect 8220 1936 8284 2000
rect 13740 1936 13804 2000
rect 13820 1936 13884 2000
rect 13900 1936 13964 2000
rect 13980 1936 14044 2000
rect 14060 1936 14124 2000
rect 14140 1936 14204 2000
rect 14220 1936 14284 2000
rect 19740 1936 19804 2000
rect 19820 1936 19884 2000
rect 19900 1936 19964 2000
rect 19980 1936 20044 2000
rect 20060 1936 20124 2000
rect 20140 1936 20204 2000
rect 20220 1936 20284 2000
rect 25740 1936 25804 2000
rect 25820 1936 25884 2000
rect 25900 1936 25964 2000
rect 25980 1936 26044 2000
rect 26060 1936 26124 2000
rect 26140 1936 26204 2000
rect 26220 1936 26284 2000
rect 31740 1936 31804 2000
rect 31820 1996 31884 2000
rect 31900 1996 31964 2000
rect 31980 1996 32044 2000
rect 32060 1996 32124 2000
rect 32140 1996 32204 2000
rect 31820 1940 31864 1996
rect 31864 1940 31884 1996
rect 31900 1940 31920 1996
rect 31920 1940 31944 1996
rect 31944 1940 31964 1996
rect 31980 1940 32000 1996
rect 32000 1940 32024 1996
rect 32024 1940 32044 1996
rect 32060 1940 32080 1996
rect 32080 1940 32104 1996
rect 32104 1940 32124 1996
rect 32140 1940 32160 1996
rect 32160 1940 32204 1996
rect 31820 1936 31884 1940
rect 31900 1936 31964 1940
rect 31980 1936 32044 1940
rect 32060 1936 32124 1940
rect 32140 1936 32204 1940
rect 32220 1936 32284 2000
rect 37740 1936 37804 2000
rect 37820 1936 37884 2000
rect 37900 1936 37964 2000
rect 37980 1936 38044 2000
rect 38060 1936 38124 2000
rect 38140 1936 38204 2000
rect 38220 1936 38284 2000
rect 43740 1936 43804 2000
rect 43820 1936 43884 2000
rect 43900 1936 43964 2000
rect 43980 1936 44044 2000
rect 44060 1936 44124 2000
rect 44140 1936 44204 2000
rect 44220 1936 44284 2000
rect 49740 1936 49804 2000
rect 49820 1936 49884 2000
rect 49900 1936 49964 2000
rect 49980 1936 50044 2000
rect 50060 1936 50124 2000
rect 50140 1936 50204 2000
rect 50220 1936 50284 2000
rect 55740 1936 55804 2000
rect 55820 1936 55884 2000
rect 55900 1936 55964 2000
rect 55980 1936 56044 2000
rect 56060 1936 56124 2000
rect 56140 1936 56204 2000
rect 56220 1936 56284 2000
rect 61740 1936 61804 2000
rect 61820 1996 61884 2000
rect 61900 1996 61964 2000
rect 61980 1996 62044 2000
rect 62060 1996 62124 2000
rect 62140 1996 62204 2000
rect 61820 1940 61864 1996
rect 61864 1940 61884 1996
rect 61900 1940 61920 1996
rect 61920 1940 61944 1996
rect 61944 1940 61964 1996
rect 61980 1940 62000 1996
rect 62000 1940 62024 1996
rect 62024 1940 62044 1996
rect 62060 1940 62080 1996
rect 62080 1940 62104 1996
rect 62104 1940 62124 1996
rect 62140 1940 62160 1996
rect 62160 1940 62204 1996
rect 61820 1936 61884 1940
rect 61900 1936 61964 1940
rect 61980 1936 62044 1940
rect 62060 1936 62124 1940
rect 62140 1936 62204 1940
rect 62220 1936 62284 2000
rect 67740 1936 67804 2000
rect 67820 1936 67884 2000
rect 67900 1936 67964 2000
rect 67980 1936 68044 2000
rect 68060 1936 68124 2000
rect 68140 1936 68204 2000
rect 68220 1936 68284 2000
rect 73740 1936 73804 2000
rect 73820 1936 73884 2000
rect 73900 1936 73964 2000
rect 73980 1936 74044 2000
rect 74060 1936 74124 2000
rect 74140 1936 74204 2000
rect 74220 1936 74284 2000
<< metal4 >>
rect 1702 82240 2322 87000
rect 1702 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82176 2220 82240
rect 2284 82176 2322 82240
rect 1702 82160 2322 82176
rect 1702 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82096 2220 82160
rect 2284 82096 2322 82160
rect 1702 82080 2322 82096
rect 1702 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82016 2220 82080
rect 2284 82016 2322 82080
rect 1702 82000 2322 82016
rect 1702 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81936 2220 82000
rect 2284 81936 2322 82000
rect 1702 72240 2322 81936
rect 1702 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72176 2220 72240
rect 2284 72176 2322 72240
rect 1702 72160 2322 72176
rect 1702 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72096 2220 72160
rect 2284 72096 2322 72160
rect 1702 72080 2322 72096
rect 1702 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72016 2220 72080
rect 2284 72016 2322 72080
rect 1702 72000 2322 72016
rect 1702 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71936 2220 72000
rect 2284 71936 2322 72000
rect 1702 62240 2322 71936
rect 1702 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62176 2220 62240
rect 2284 62176 2322 62240
rect 1702 62160 2322 62176
rect 1702 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62096 2220 62160
rect 2284 62096 2322 62160
rect 1702 62080 2322 62096
rect 1702 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62016 2220 62080
rect 2284 62016 2322 62080
rect 1702 62000 2322 62016
rect 1702 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61936 2220 62000
rect 2284 61936 2322 62000
rect 1702 52240 2322 61936
rect 1702 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52176 2220 52240
rect 2284 52176 2322 52240
rect 1702 52160 2322 52176
rect 1702 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52096 2220 52160
rect 2284 52096 2322 52160
rect 1702 52080 2322 52096
rect 1702 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52016 2220 52080
rect 2284 52016 2322 52080
rect 1702 52000 2322 52016
rect 1702 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51936 2220 52000
rect 2284 51936 2322 52000
rect 1702 42240 2322 51936
rect 1702 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42176 2220 42240
rect 2284 42176 2322 42240
rect 1702 42160 2322 42176
rect 1702 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42096 2220 42160
rect 2284 42096 2322 42160
rect 1702 42080 2322 42096
rect 1702 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42016 2220 42080
rect 2284 42016 2322 42080
rect 1702 42000 2322 42016
rect 1702 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41936 2220 42000
rect 2284 41936 2322 42000
rect 1702 32240 2322 41936
rect 1702 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32176 2220 32240
rect 2284 32176 2322 32240
rect 1702 32160 2322 32176
rect 1702 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32096 2220 32160
rect 2284 32096 2322 32160
rect 1702 32080 2322 32096
rect 1702 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32016 2220 32080
rect 2284 32016 2322 32080
rect 1702 32000 2322 32016
rect 1702 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31936 2220 32000
rect 2284 31936 2322 32000
rect 1702 22240 2322 31936
rect 1702 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22176 2220 22240
rect 2284 22176 2322 22240
rect 1702 22160 2322 22176
rect 1702 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22096 2220 22160
rect 2284 22096 2322 22160
rect 1702 22080 2322 22096
rect 1702 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22016 2220 22080
rect 2284 22016 2322 22080
rect 1702 22000 2322 22016
rect 1702 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21936 2220 22000
rect 2284 21936 2322 22000
rect 1702 12240 2322 21936
rect 1702 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12176 2220 12240
rect 2284 12176 2322 12240
rect 1702 12160 2322 12176
rect 1702 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12096 2220 12160
rect 2284 12096 2322 12160
rect 1702 12080 2322 12096
rect 1702 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12016 2220 12080
rect 2284 12016 2322 12080
rect 1702 12000 2322 12016
rect 1702 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2220 12000
rect 2284 11936 2322 12000
rect 1702 2240 2322 11936
rect 1702 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2176 1900 2240
rect 1964 2176 1980 2240
rect 2044 2176 2060 2240
rect 2124 2176 2140 2240
rect 2204 2176 2220 2240
rect 2284 2176 2322 2240
rect 1702 2160 2322 2176
rect 1702 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2096 1900 2160
rect 1964 2096 1980 2160
rect 2044 2096 2060 2160
rect 2124 2096 2140 2160
rect 2204 2096 2220 2160
rect 2284 2096 2322 2160
rect 1702 2080 2322 2096
rect 1702 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2016 1900 2080
rect 1964 2016 1980 2080
rect 2044 2016 2060 2080
rect 2124 2016 2140 2080
rect 2204 2016 2220 2080
rect 2284 2016 2322 2080
rect 1702 2000 2322 2016
rect 1702 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1936 1900 2000
rect 1964 1936 1980 2000
rect 2044 1936 2060 2000
rect 2124 1936 2140 2000
rect 2204 1936 2220 2000
rect 2284 1936 2322 2000
rect 1702 0 2322 1936
rect 4702 84592 5322 87000
rect 4702 84528 4740 84592
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84528 5322 84592
rect 4702 84512 5322 84528
rect 4702 84448 4740 84512
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84448 5322 84512
rect 4702 84432 5322 84448
rect 4702 84368 4740 84432
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84368 5322 84432
rect 4702 84352 5322 84368
rect 4702 84288 4740 84352
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84288 5322 84352
rect 4702 74592 5322 84288
rect 4702 74528 4740 74592
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74528 5322 74592
rect 4702 74512 5322 74528
rect 4702 74448 4740 74512
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74448 5322 74512
rect 4702 74432 5322 74448
rect 4702 74368 4740 74432
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74368 5322 74432
rect 4702 74352 5322 74368
rect 4702 74288 4740 74352
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74288 5322 74352
rect 4702 64592 5322 74288
rect 4702 64528 4740 64592
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64528 5322 64592
rect 4702 64512 5322 64528
rect 4702 64448 4740 64512
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64448 5322 64512
rect 4702 64432 5322 64448
rect 4702 64368 4740 64432
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64368 5322 64432
rect 4702 64352 5322 64368
rect 4702 64288 4740 64352
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64288 5322 64352
rect 4702 54592 5322 64288
rect 4702 54528 4740 54592
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54528 5322 54592
rect 4702 54512 5322 54528
rect 4702 54448 4740 54512
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54448 5322 54512
rect 4702 54432 5322 54448
rect 4702 54368 4740 54432
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54368 5322 54432
rect 4702 54352 5322 54368
rect 4702 54288 4740 54352
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54288 5322 54352
rect 4702 44592 5322 54288
rect 4702 44528 4740 44592
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44528 5322 44592
rect 4702 44512 5322 44528
rect 4702 44448 4740 44512
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44448 5322 44512
rect 4702 44432 5322 44448
rect 4702 44368 4740 44432
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44368 5322 44432
rect 4702 44352 5322 44368
rect 4702 44288 4740 44352
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44288 5322 44352
rect 4702 34592 5322 44288
rect 4702 34528 4740 34592
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34528 5322 34592
rect 4702 34512 5322 34528
rect 4702 34448 4740 34512
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34448 5322 34512
rect 4702 34432 5322 34448
rect 4702 34368 4740 34432
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34368 5322 34432
rect 4702 34352 5322 34368
rect 4702 34288 4740 34352
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34288 5322 34352
rect 4702 24592 5322 34288
rect 4702 24528 4740 24592
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24528 5322 24592
rect 4702 24512 5322 24528
rect 4702 24448 4740 24512
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24448 5322 24512
rect 4702 24432 5322 24448
rect 4702 24368 4740 24432
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24368 5322 24432
rect 4702 24352 5322 24368
rect 4702 24288 4740 24352
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24288 5322 24352
rect 4702 14592 5322 24288
rect 4702 14528 4740 14592
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14528 5322 14592
rect 4702 14512 5322 14528
rect 4702 14448 4740 14512
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14448 5322 14512
rect 4702 14432 5322 14448
rect 4702 14368 4740 14432
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14368 5322 14432
rect 4702 14352 5322 14368
rect 4702 14288 4740 14352
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14288 5322 14352
rect 4702 4592 5322 14288
rect 4702 4528 4740 4592
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 5322 4592
rect 4702 4512 5322 4528
rect 4702 4448 4740 4512
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 5322 4512
rect 4702 4432 5322 4448
rect 4702 4368 4740 4432
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 5322 4432
rect 4702 4352 5322 4368
rect 4702 4288 4740 4352
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 5322 4352
rect 4702 0 5322 4288
rect 7702 82240 8322 87000
rect 7702 82176 7740 82240
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82176 8322 82240
rect 7702 82160 8322 82176
rect 7702 82096 7740 82160
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82096 8322 82160
rect 7702 82080 8322 82096
rect 7702 82016 7740 82080
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82016 8322 82080
rect 7702 82000 8322 82016
rect 7702 81936 7740 82000
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81936 8322 82000
rect 7702 72240 8322 81936
rect 7702 72176 7740 72240
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72176 8322 72240
rect 7702 72160 8322 72176
rect 7702 72096 7740 72160
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72096 8322 72160
rect 7702 72080 8322 72096
rect 7702 72016 7740 72080
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72016 8322 72080
rect 7702 72000 8322 72016
rect 7702 71936 7740 72000
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71936 8322 72000
rect 7702 62240 8322 71936
rect 7702 62176 7740 62240
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62176 8322 62240
rect 7702 62160 8322 62176
rect 7702 62096 7740 62160
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62096 8322 62160
rect 7702 62080 8322 62096
rect 7702 62016 7740 62080
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62016 8322 62080
rect 7702 62000 8322 62016
rect 7702 61936 7740 62000
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61936 8322 62000
rect 7702 52240 8322 61936
rect 7702 52176 7740 52240
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52176 8322 52240
rect 7702 52160 8322 52176
rect 7702 52096 7740 52160
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52096 8322 52160
rect 7702 52080 8322 52096
rect 7702 52016 7740 52080
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52016 8322 52080
rect 7702 52000 8322 52016
rect 7702 51936 7740 52000
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51936 8322 52000
rect 7702 42240 8322 51936
rect 7702 42176 7740 42240
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42176 8322 42240
rect 7702 42160 8322 42176
rect 7702 42096 7740 42160
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42096 8322 42160
rect 7702 42080 8322 42096
rect 7702 42016 7740 42080
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42016 8322 42080
rect 7702 42000 8322 42016
rect 7702 41936 7740 42000
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41936 8322 42000
rect 7702 32240 8322 41936
rect 7702 32176 7740 32240
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32176 8322 32240
rect 7702 32160 8322 32176
rect 7702 32096 7740 32160
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32096 8322 32160
rect 7702 32080 8322 32096
rect 7702 32016 7740 32080
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32016 8322 32080
rect 7702 32000 8322 32016
rect 7702 31936 7740 32000
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31936 8322 32000
rect 7702 22240 8322 31936
rect 7702 22176 7740 22240
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22176 8322 22240
rect 7702 22160 8322 22176
rect 7702 22096 7740 22160
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22096 8322 22160
rect 7702 22080 8322 22096
rect 7702 22016 7740 22080
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22016 8322 22080
rect 7702 22000 8322 22016
rect 7702 21936 7740 22000
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21936 8322 22000
rect 7702 12240 8322 21936
rect 7702 12176 7740 12240
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12176 8322 12240
rect 7702 12160 8322 12176
rect 7702 12096 7740 12160
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12096 8322 12160
rect 7702 12080 8322 12096
rect 7702 12016 7740 12080
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12016 8322 12080
rect 7702 12000 8322 12016
rect 7702 11936 7740 12000
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11936 8322 12000
rect 7702 2240 8322 11936
rect 7702 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2176 8322 2240
rect 7702 2160 8322 2176
rect 7702 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2096 8322 2160
rect 7702 2080 8322 2096
rect 7702 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2016 8322 2080
rect 7702 2000 8322 2016
rect 7702 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1936 8322 2000
rect 7702 0 8322 1936
rect 10702 84592 11322 87000
rect 10702 84528 10740 84592
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84528 11322 84592
rect 10702 84512 11322 84528
rect 10702 84448 10740 84512
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84448 11322 84512
rect 10702 84432 11322 84448
rect 10702 84368 10740 84432
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84368 11322 84432
rect 10702 84352 11322 84368
rect 10702 84288 10740 84352
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84288 11322 84352
rect 10702 74592 11322 84288
rect 10702 74528 10740 74592
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74528 11322 74592
rect 10702 74512 11322 74528
rect 10702 74448 10740 74512
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74448 11322 74512
rect 10702 74432 11322 74448
rect 10702 74368 10740 74432
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74368 11322 74432
rect 10702 74352 11322 74368
rect 10702 74288 10740 74352
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74288 11322 74352
rect 10702 64592 11322 74288
rect 10702 64528 10740 64592
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64528 11322 64592
rect 10702 64512 11322 64528
rect 10702 64448 10740 64512
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64448 11322 64512
rect 10702 64432 11322 64448
rect 10702 64368 10740 64432
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64368 11322 64432
rect 10702 64352 11322 64368
rect 10702 64288 10740 64352
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64288 11322 64352
rect 10702 54592 11322 64288
rect 10702 54528 10740 54592
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54528 11322 54592
rect 10702 54512 11322 54528
rect 10702 54448 10740 54512
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54448 11322 54512
rect 10702 54432 11322 54448
rect 10702 54368 10740 54432
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54368 11322 54432
rect 10702 54352 11322 54368
rect 10702 54288 10740 54352
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54288 11322 54352
rect 10702 44592 11322 54288
rect 10702 44528 10740 44592
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44528 11322 44592
rect 10702 44512 11322 44528
rect 10702 44448 10740 44512
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44448 11322 44512
rect 10702 44432 11322 44448
rect 10702 44368 10740 44432
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44368 11322 44432
rect 10702 44352 11322 44368
rect 10702 44288 10740 44352
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44288 11322 44352
rect 10702 34592 11322 44288
rect 10702 34528 10740 34592
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34528 11322 34592
rect 10702 34512 11322 34528
rect 10702 34448 10740 34512
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34448 11322 34512
rect 10702 34432 11322 34448
rect 10702 34368 10740 34432
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34368 11322 34432
rect 10702 34352 11322 34368
rect 10702 34288 10740 34352
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34288 11322 34352
rect 10702 24592 11322 34288
rect 10702 24528 10740 24592
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24528 11322 24592
rect 10702 24512 11322 24528
rect 10702 24448 10740 24512
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24448 11322 24512
rect 10702 24432 11322 24448
rect 10702 24368 10740 24432
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24368 11322 24432
rect 10702 24352 11322 24368
rect 10702 24288 10740 24352
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24288 11322 24352
rect 10702 14592 11322 24288
rect 10702 14528 10740 14592
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14528 11322 14592
rect 10702 14512 11322 14528
rect 10702 14448 10740 14512
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14448 11322 14512
rect 10702 14432 11322 14448
rect 10702 14368 10740 14432
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14368 11322 14432
rect 10702 14352 11322 14368
rect 10702 14288 10740 14352
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14288 11322 14352
rect 10702 4592 11322 14288
rect 10702 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4528 11322 4592
rect 10702 4512 11322 4528
rect 10702 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4448 11322 4512
rect 10702 4432 11322 4448
rect 10702 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4368 11322 4432
rect 10702 4352 11322 4368
rect 10702 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4288 11322 4352
rect 10702 0 11322 4288
rect 13702 82240 14322 87000
rect 13702 82176 13740 82240
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82176 14220 82240
rect 14284 82176 14322 82240
rect 13702 82160 14322 82176
rect 13702 82096 13740 82160
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82096 14220 82160
rect 14284 82096 14322 82160
rect 13702 82080 14322 82096
rect 13702 82016 13740 82080
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82016 14220 82080
rect 14284 82016 14322 82080
rect 13702 82000 14322 82016
rect 13702 81936 13740 82000
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81936 14220 82000
rect 14284 81936 14322 82000
rect 13702 72240 14322 81936
rect 13702 72176 13740 72240
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72176 14220 72240
rect 14284 72176 14322 72240
rect 13702 72160 14322 72176
rect 13702 72096 13740 72160
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72096 14220 72160
rect 14284 72096 14322 72160
rect 13702 72080 14322 72096
rect 13702 72016 13740 72080
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72016 14220 72080
rect 14284 72016 14322 72080
rect 13702 72000 14322 72016
rect 13702 71936 13740 72000
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71936 14220 72000
rect 14284 71936 14322 72000
rect 13702 62240 14322 71936
rect 13702 62176 13740 62240
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62176 14220 62240
rect 14284 62176 14322 62240
rect 13702 62160 14322 62176
rect 13702 62096 13740 62160
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62096 14220 62160
rect 14284 62096 14322 62160
rect 13702 62080 14322 62096
rect 13702 62016 13740 62080
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62016 14220 62080
rect 14284 62016 14322 62080
rect 13702 62000 14322 62016
rect 13702 61936 13740 62000
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61936 14220 62000
rect 14284 61936 14322 62000
rect 13702 52240 14322 61936
rect 13702 52176 13740 52240
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52176 14220 52240
rect 14284 52176 14322 52240
rect 13702 52160 14322 52176
rect 13702 52096 13740 52160
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52096 14220 52160
rect 14284 52096 14322 52160
rect 13702 52080 14322 52096
rect 13702 52016 13740 52080
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52016 14220 52080
rect 14284 52016 14322 52080
rect 13702 52000 14322 52016
rect 13702 51936 13740 52000
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51936 14220 52000
rect 14284 51936 14322 52000
rect 13702 42240 14322 51936
rect 13702 42176 13740 42240
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42176 14220 42240
rect 14284 42176 14322 42240
rect 13702 42160 14322 42176
rect 13702 42096 13740 42160
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42096 14220 42160
rect 14284 42096 14322 42160
rect 13702 42080 14322 42096
rect 13702 42016 13740 42080
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42016 14220 42080
rect 14284 42016 14322 42080
rect 13702 42000 14322 42016
rect 13702 41936 13740 42000
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41936 14220 42000
rect 14284 41936 14322 42000
rect 13702 32240 14322 41936
rect 13702 32176 13740 32240
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32176 14220 32240
rect 14284 32176 14322 32240
rect 13702 32160 14322 32176
rect 13702 32096 13740 32160
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32096 14220 32160
rect 14284 32096 14322 32160
rect 13702 32080 14322 32096
rect 13702 32016 13740 32080
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32016 14220 32080
rect 14284 32016 14322 32080
rect 13702 32000 14322 32016
rect 13702 31936 13740 32000
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31936 14220 32000
rect 14284 31936 14322 32000
rect 13702 22240 14322 31936
rect 13702 22176 13740 22240
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22176 14220 22240
rect 14284 22176 14322 22240
rect 13702 22160 14322 22176
rect 13702 22096 13740 22160
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22096 14220 22160
rect 14284 22096 14322 22160
rect 13702 22080 14322 22096
rect 13702 22016 13740 22080
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22016 14220 22080
rect 14284 22016 14322 22080
rect 13702 22000 14322 22016
rect 13702 21936 13740 22000
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21936 14220 22000
rect 14284 21936 14322 22000
rect 13702 12240 14322 21936
rect 13702 12176 13740 12240
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12176 14220 12240
rect 14284 12176 14322 12240
rect 13702 12160 14322 12176
rect 13702 12096 13740 12160
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12096 14220 12160
rect 14284 12096 14322 12160
rect 13702 12080 14322 12096
rect 13702 12016 13740 12080
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12016 14220 12080
rect 14284 12016 14322 12080
rect 13702 12000 14322 12016
rect 13702 11936 13740 12000
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11936 14220 12000
rect 14284 11936 14322 12000
rect 13702 2240 14322 11936
rect 13702 2176 13740 2240
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 14322 2240
rect 13702 2160 14322 2176
rect 13702 2096 13740 2160
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 14322 2160
rect 13702 2080 14322 2096
rect 13702 2016 13740 2080
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 14322 2080
rect 13702 2000 14322 2016
rect 13702 1936 13740 2000
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 14322 2000
rect 13702 0 14322 1936
rect 16702 84592 17322 87000
rect 16702 84528 16740 84592
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84528 17140 84592
rect 17204 84528 17220 84592
rect 17284 84528 17322 84592
rect 16702 84512 17322 84528
rect 16702 84448 16740 84512
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84448 17140 84512
rect 17204 84448 17220 84512
rect 17284 84448 17322 84512
rect 16702 84432 17322 84448
rect 16702 84368 16740 84432
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84368 17140 84432
rect 17204 84368 17220 84432
rect 17284 84368 17322 84432
rect 16702 84352 17322 84368
rect 16702 84288 16740 84352
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84288 17140 84352
rect 17204 84288 17220 84352
rect 17284 84288 17322 84352
rect 16702 74592 17322 84288
rect 16702 74528 16740 74592
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74528 17140 74592
rect 17204 74528 17220 74592
rect 17284 74528 17322 74592
rect 16702 74512 17322 74528
rect 16702 74448 16740 74512
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74448 17140 74512
rect 17204 74448 17220 74512
rect 17284 74448 17322 74512
rect 16702 74432 17322 74448
rect 16702 74368 16740 74432
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74368 17140 74432
rect 17204 74368 17220 74432
rect 17284 74368 17322 74432
rect 16702 74352 17322 74368
rect 16702 74288 16740 74352
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74288 17140 74352
rect 17204 74288 17220 74352
rect 17284 74288 17322 74352
rect 16702 64592 17322 74288
rect 16702 64528 16740 64592
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64528 17140 64592
rect 17204 64528 17220 64592
rect 17284 64528 17322 64592
rect 16702 64512 17322 64528
rect 16702 64448 16740 64512
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64448 17140 64512
rect 17204 64448 17220 64512
rect 17284 64448 17322 64512
rect 16702 64432 17322 64448
rect 16702 64368 16740 64432
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64368 17140 64432
rect 17204 64368 17220 64432
rect 17284 64368 17322 64432
rect 16702 64352 17322 64368
rect 16702 64288 16740 64352
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64288 17140 64352
rect 17204 64288 17220 64352
rect 17284 64288 17322 64352
rect 16702 54592 17322 64288
rect 16702 54528 16740 54592
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54528 17140 54592
rect 17204 54528 17220 54592
rect 17284 54528 17322 54592
rect 16702 54512 17322 54528
rect 16702 54448 16740 54512
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54448 17140 54512
rect 17204 54448 17220 54512
rect 17284 54448 17322 54512
rect 16702 54432 17322 54448
rect 16702 54368 16740 54432
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54368 17140 54432
rect 17204 54368 17220 54432
rect 17284 54368 17322 54432
rect 16702 54352 17322 54368
rect 16702 54288 16740 54352
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54288 17140 54352
rect 17204 54288 17220 54352
rect 17284 54288 17322 54352
rect 16702 44592 17322 54288
rect 16702 44528 16740 44592
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44528 17140 44592
rect 17204 44528 17220 44592
rect 17284 44528 17322 44592
rect 16702 44512 17322 44528
rect 16702 44448 16740 44512
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44448 17140 44512
rect 17204 44448 17220 44512
rect 17284 44448 17322 44512
rect 16702 44432 17322 44448
rect 16702 44368 16740 44432
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44368 17140 44432
rect 17204 44368 17220 44432
rect 17284 44368 17322 44432
rect 16702 44352 17322 44368
rect 16702 44288 16740 44352
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44288 17140 44352
rect 17204 44288 17220 44352
rect 17284 44288 17322 44352
rect 16702 34592 17322 44288
rect 16702 34528 16740 34592
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34528 17140 34592
rect 17204 34528 17220 34592
rect 17284 34528 17322 34592
rect 16702 34512 17322 34528
rect 16702 34448 16740 34512
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34448 17140 34512
rect 17204 34448 17220 34512
rect 17284 34448 17322 34512
rect 16702 34432 17322 34448
rect 16702 34368 16740 34432
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34368 17140 34432
rect 17204 34368 17220 34432
rect 17284 34368 17322 34432
rect 16702 34352 17322 34368
rect 16702 34288 16740 34352
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34288 17140 34352
rect 17204 34288 17220 34352
rect 17284 34288 17322 34352
rect 16702 24592 17322 34288
rect 16702 24528 16740 24592
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24528 17140 24592
rect 17204 24528 17220 24592
rect 17284 24528 17322 24592
rect 16702 24512 17322 24528
rect 16702 24448 16740 24512
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24448 17140 24512
rect 17204 24448 17220 24512
rect 17284 24448 17322 24512
rect 16702 24432 17322 24448
rect 16702 24368 16740 24432
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24368 17140 24432
rect 17204 24368 17220 24432
rect 17284 24368 17322 24432
rect 16702 24352 17322 24368
rect 16702 24288 16740 24352
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24288 17140 24352
rect 17204 24288 17220 24352
rect 17284 24288 17322 24352
rect 16702 14592 17322 24288
rect 16702 14528 16740 14592
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14528 17140 14592
rect 17204 14528 17220 14592
rect 17284 14528 17322 14592
rect 16702 14512 17322 14528
rect 16702 14448 16740 14512
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14448 17140 14512
rect 17204 14448 17220 14512
rect 17284 14448 17322 14512
rect 16702 14432 17322 14448
rect 16702 14368 16740 14432
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14368 17140 14432
rect 17204 14368 17220 14432
rect 17284 14368 17322 14432
rect 16702 14352 17322 14368
rect 16702 14288 16740 14352
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14288 17140 14352
rect 17204 14288 17220 14352
rect 17284 14288 17322 14352
rect 16702 4592 17322 14288
rect 16702 4528 16740 4592
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 17322 4592
rect 16702 4512 17322 4528
rect 16702 4448 16740 4512
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 17322 4512
rect 16702 4432 17322 4448
rect 16702 4368 16740 4432
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 17322 4432
rect 16702 4352 17322 4368
rect 16702 4288 16740 4352
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 17322 4352
rect 16702 0 17322 4288
rect 19702 82240 20322 87000
rect 19702 82176 19740 82240
rect 19804 82176 19820 82240
rect 19884 82176 19900 82240
rect 19964 82176 19980 82240
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82176 20322 82240
rect 19702 82160 20322 82176
rect 19702 82096 19740 82160
rect 19804 82096 19820 82160
rect 19884 82096 19900 82160
rect 19964 82096 19980 82160
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82096 20322 82160
rect 19702 82080 20322 82096
rect 19702 82016 19740 82080
rect 19804 82016 19820 82080
rect 19884 82016 19900 82080
rect 19964 82016 19980 82080
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82016 20322 82080
rect 19702 82000 20322 82016
rect 19702 81936 19740 82000
rect 19804 81936 19820 82000
rect 19884 81936 19900 82000
rect 19964 81936 19980 82000
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81936 20322 82000
rect 19702 72240 20322 81936
rect 19702 72176 19740 72240
rect 19804 72176 19820 72240
rect 19884 72176 19900 72240
rect 19964 72176 19980 72240
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72176 20322 72240
rect 19702 72160 20322 72176
rect 19702 72096 19740 72160
rect 19804 72096 19820 72160
rect 19884 72096 19900 72160
rect 19964 72096 19980 72160
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72096 20322 72160
rect 19702 72080 20322 72096
rect 19702 72016 19740 72080
rect 19804 72016 19820 72080
rect 19884 72016 19900 72080
rect 19964 72016 19980 72080
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72016 20322 72080
rect 19702 72000 20322 72016
rect 19702 71936 19740 72000
rect 19804 71936 19820 72000
rect 19884 71936 19900 72000
rect 19964 71936 19980 72000
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71936 20322 72000
rect 19702 62240 20322 71936
rect 19702 62176 19740 62240
rect 19804 62176 19820 62240
rect 19884 62176 19900 62240
rect 19964 62176 19980 62240
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62176 20322 62240
rect 19702 62160 20322 62176
rect 19702 62096 19740 62160
rect 19804 62096 19820 62160
rect 19884 62096 19900 62160
rect 19964 62096 19980 62160
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62096 20322 62160
rect 19702 62080 20322 62096
rect 19702 62016 19740 62080
rect 19804 62016 19820 62080
rect 19884 62016 19900 62080
rect 19964 62016 19980 62080
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62016 20322 62080
rect 19702 62000 20322 62016
rect 19702 61936 19740 62000
rect 19804 61936 19820 62000
rect 19884 61936 19900 62000
rect 19964 61936 19980 62000
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61936 20322 62000
rect 19702 52240 20322 61936
rect 19702 52176 19740 52240
rect 19804 52176 19820 52240
rect 19884 52176 19900 52240
rect 19964 52176 19980 52240
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52176 20322 52240
rect 19702 52160 20322 52176
rect 19702 52096 19740 52160
rect 19804 52096 19820 52160
rect 19884 52096 19900 52160
rect 19964 52096 19980 52160
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52096 20322 52160
rect 19702 52080 20322 52096
rect 19702 52016 19740 52080
rect 19804 52016 19820 52080
rect 19884 52016 19900 52080
rect 19964 52016 19980 52080
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52016 20322 52080
rect 19702 52000 20322 52016
rect 19702 51936 19740 52000
rect 19804 51936 19820 52000
rect 19884 51936 19900 52000
rect 19964 51936 19980 52000
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51936 20322 52000
rect 19702 42240 20322 51936
rect 19702 42176 19740 42240
rect 19804 42176 19820 42240
rect 19884 42176 19900 42240
rect 19964 42176 19980 42240
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42176 20322 42240
rect 19702 42160 20322 42176
rect 19702 42096 19740 42160
rect 19804 42096 19820 42160
rect 19884 42096 19900 42160
rect 19964 42096 19980 42160
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42096 20322 42160
rect 19702 42080 20322 42096
rect 19702 42016 19740 42080
rect 19804 42016 19820 42080
rect 19884 42016 19900 42080
rect 19964 42016 19980 42080
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42016 20322 42080
rect 19702 42000 20322 42016
rect 19702 41936 19740 42000
rect 19804 41936 19820 42000
rect 19884 41936 19900 42000
rect 19964 41936 19980 42000
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41936 20322 42000
rect 19702 32240 20322 41936
rect 19702 32176 19740 32240
rect 19804 32176 19820 32240
rect 19884 32176 19900 32240
rect 19964 32176 19980 32240
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32176 20322 32240
rect 19702 32160 20322 32176
rect 19702 32096 19740 32160
rect 19804 32096 19820 32160
rect 19884 32096 19900 32160
rect 19964 32096 19980 32160
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32096 20322 32160
rect 19702 32080 20322 32096
rect 19702 32016 19740 32080
rect 19804 32016 19820 32080
rect 19884 32016 19900 32080
rect 19964 32016 19980 32080
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32016 20322 32080
rect 19702 32000 20322 32016
rect 19702 31936 19740 32000
rect 19804 31936 19820 32000
rect 19884 31936 19900 32000
rect 19964 31936 19980 32000
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31936 20322 32000
rect 19702 22240 20322 31936
rect 19702 22176 19740 22240
rect 19804 22176 19820 22240
rect 19884 22176 19900 22240
rect 19964 22176 19980 22240
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22176 20322 22240
rect 19702 22160 20322 22176
rect 19702 22096 19740 22160
rect 19804 22096 19820 22160
rect 19884 22096 19900 22160
rect 19964 22096 19980 22160
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22096 20322 22160
rect 19702 22080 20322 22096
rect 19702 22016 19740 22080
rect 19804 22016 19820 22080
rect 19884 22016 19900 22080
rect 19964 22016 19980 22080
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22016 20322 22080
rect 19702 22000 20322 22016
rect 19702 21936 19740 22000
rect 19804 21936 19820 22000
rect 19884 21936 19900 22000
rect 19964 21936 19980 22000
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21936 20322 22000
rect 19702 12240 20322 21936
rect 19702 12176 19740 12240
rect 19804 12176 19820 12240
rect 19884 12176 19900 12240
rect 19964 12176 19980 12240
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12176 20322 12240
rect 19702 12160 20322 12176
rect 19702 12096 19740 12160
rect 19804 12096 19820 12160
rect 19884 12096 19900 12160
rect 19964 12096 19980 12160
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12096 20322 12160
rect 19702 12080 20322 12096
rect 19702 12016 19740 12080
rect 19804 12016 19820 12080
rect 19884 12016 19900 12080
rect 19964 12016 19980 12080
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12016 20322 12080
rect 19702 12000 20322 12016
rect 19702 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11936 20322 12000
rect 19702 2240 20322 11936
rect 19702 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2176 20322 2240
rect 19702 2160 20322 2176
rect 19702 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2096 20322 2160
rect 19702 2080 20322 2096
rect 19702 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2016 20322 2080
rect 19702 2000 20322 2016
rect 19702 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1936 20322 2000
rect 19702 0 20322 1936
rect 22702 84592 23322 87000
rect 22702 84528 22740 84592
rect 22804 84528 22820 84592
rect 22884 84528 22900 84592
rect 22964 84528 22980 84592
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84528 23322 84592
rect 22702 84512 23322 84528
rect 22702 84448 22740 84512
rect 22804 84448 22820 84512
rect 22884 84448 22900 84512
rect 22964 84448 22980 84512
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84448 23322 84512
rect 22702 84432 23322 84448
rect 22702 84368 22740 84432
rect 22804 84368 22820 84432
rect 22884 84368 22900 84432
rect 22964 84368 22980 84432
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84368 23322 84432
rect 22702 84352 23322 84368
rect 22702 84288 22740 84352
rect 22804 84288 22820 84352
rect 22884 84288 22900 84352
rect 22964 84288 22980 84352
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84288 23322 84352
rect 22702 74592 23322 84288
rect 22702 74528 22740 74592
rect 22804 74528 22820 74592
rect 22884 74528 22900 74592
rect 22964 74528 22980 74592
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74528 23322 74592
rect 22702 74512 23322 74528
rect 22702 74448 22740 74512
rect 22804 74448 22820 74512
rect 22884 74448 22900 74512
rect 22964 74448 22980 74512
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74448 23322 74512
rect 22702 74432 23322 74448
rect 22702 74368 22740 74432
rect 22804 74368 22820 74432
rect 22884 74368 22900 74432
rect 22964 74368 22980 74432
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74368 23322 74432
rect 22702 74352 23322 74368
rect 22702 74288 22740 74352
rect 22804 74288 22820 74352
rect 22884 74288 22900 74352
rect 22964 74288 22980 74352
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74288 23322 74352
rect 22702 64592 23322 74288
rect 22702 64528 22740 64592
rect 22804 64528 22820 64592
rect 22884 64528 22900 64592
rect 22964 64528 22980 64592
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64528 23322 64592
rect 22702 64512 23322 64528
rect 22702 64448 22740 64512
rect 22804 64448 22820 64512
rect 22884 64448 22900 64512
rect 22964 64448 22980 64512
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64448 23322 64512
rect 22702 64432 23322 64448
rect 22702 64368 22740 64432
rect 22804 64368 22820 64432
rect 22884 64368 22900 64432
rect 22964 64368 22980 64432
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64368 23322 64432
rect 22702 64352 23322 64368
rect 22702 64288 22740 64352
rect 22804 64288 22820 64352
rect 22884 64288 22900 64352
rect 22964 64288 22980 64352
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64288 23322 64352
rect 22702 54592 23322 64288
rect 22702 54528 22740 54592
rect 22804 54528 22820 54592
rect 22884 54528 22900 54592
rect 22964 54528 22980 54592
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54528 23322 54592
rect 22702 54512 23322 54528
rect 22702 54448 22740 54512
rect 22804 54448 22820 54512
rect 22884 54448 22900 54512
rect 22964 54448 22980 54512
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54448 23322 54512
rect 22702 54432 23322 54448
rect 22702 54368 22740 54432
rect 22804 54368 22820 54432
rect 22884 54368 22900 54432
rect 22964 54368 22980 54432
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54368 23322 54432
rect 22702 54352 23322 54368
rect 22702 54288 22740 54352
rect 22804 54288 22820 54352
rect 22884 54288 22900 54352
rect 22964 54288 22980 54352
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54288 23322 54352
rect 22702 44592 23322 54288
rect 22702 44528 22740 44592
rect 22804 44528 22820 44592
rect 22884 44528 22900 44592
rect 22964 44528 22980 44592
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44528 23322 44592
rect 22702 44512 23322 44528
rect 22702 44448 22740 44512
rect 22804 44448 22820 44512
rect 22884 44448 22900 44512
rect 22964 44448 22980 44512
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44448 23322 44512
rect 22702 44432 23322 44448
rect 22702 44368 22740 44432
rect 22804 44368 22820 44432
rect 22884 44368 22900 44432
rect 22964 44368 22980 44432
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44368 23322 44432
rect 22702 44352 23322 44368
rect 22702 44288 22740 44352
rect 22804 44288 22820 44352
rect 22884 44288 22900 44352
rect 22964 44288 22980 44352
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44288 23322 44352
rect 22702 34592 23322 44288
rect 22702 34528 22740 34592
rect 22804 34528 22820 34592
rect 22884 34528 22900 34592
rect 22964 34528 22980 34592
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34528 23322 34592
rect 22702 34512 23322 34528
rect 22702 34448 22740 34512
rect 22804 34448 22820 34512
rect 22884 34448 22900 34512
rect 22964 34448 22980 34512
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34448 23322 34512
rect 22702 34432 23322 34448
rect 22702 34368 22740 34432
rect 22804 34368 22820 34432
rect 22884 34368 22900 34432
rect 22964 34368 22980 34432
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34368 23322 34432
rect 22702 34352 23322 34368
rect 22702 34288 22740 34352
rect 22804 34288 22820 34352
rect 22884 34288 22900 34352
rect 22964 34288 22980 34352
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34288 23322 34352
rect 22702 24592 23322 34288
rect 22702 24528 22740 24592
rect 22804 24528 22820 24592
rect 22884 24528 22900 24592
rect 22964 24528 22980 24592
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24528 23322 24592
rect 22702 24512 23322 24528
rect 22702 24448 22740 24512
rect 22804 24448 22820 24512
rect 22884 24448 22900 24512
rect 22964 24448 22980 24512
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24448 23322 24512
rect 22702 24432 23322 24448
rect 22702 24368 22740 24432
rect 22804 24368 22820 24432
rect 22884 24368 22900 24432
rect 22964 24368 22980 24432
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24368 23322 24432
rect 22702 24352 23322 24368
rect 22702 24288 22740 24352
rect 22804 24288 22820 24352
rect 22884 24288 22900 24352
rect 22964 24288 22980 24352
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24288 23322 24352
rect 22702 14592 23322 24288
rect 22702 14528 22740 14592
rect 22804 14528 22820 14592
rect 22884 14528 22900 14592
rect 22964 14528 22980 14592
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14528 23322 14592
rect 22702 14512 23322 14528
rect 22702 14448 22740 14512
rect 22804 14448 22820 14512
rect 22884 14448 22900 14512
rect 22964 14448 22980 14512
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14448 23322 14512
rect 22702 14432 23322 14448
rect 22702 14368 22740 14432
rect 22804 14368 22820 14432
rect 22884 14368 22900 14432
rect 22964 14368 22980 14432
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14368 23322 14432
rect 22702 14352 23322 14368
rect 22702 14288 22740 14352
rect 22804 14288 22820 14352
rect 22884 14288 22900 14352
rect 22964 14288 22980 14352
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14288 23322 14352
rect 22702 4592 23322 14288
rect 22702 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4528 23322 4592
rect 22702 4512 23322 4528
rect 22702 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4448 23322 4512
rect 22702 4432 23322 4448
rect 22702 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4368 23322 4432
rect 22702 4352 23322 4368
rect 22702 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4288 23322 4352
rect 22702 0 23322 4288
rect 25702 82240 26322 87000
rect 25702 82176 25740 82240
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82176 26322 82240
rect 25702 82160 26322 82176
rect 25702 82096 25740 82160
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82096 26322 82160
rect 25702 82080 26322 82096
rect 25702 82016 25740 82080
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82016 26322 82080
rect 25702 82000 26322 82016
rect 25702 81936 25740 82000
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81936 26322 82000
rect 25702 72240 26322 81936
rect 25702 72176 25740 72240
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72176 26322 72240
rect 25702 72160 26322 72176
rect 25702 72096 25740 72160
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72096 26322 72160
rect 25702 72080 26322 72096
rect 25702 72016 25740 72080
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72016 26322 72080
rect 25702 72000 26322 72016
rect 25702 71936 25740 72000
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71936 26322 72000
rect 25702 62240 26322 71936
rect 25702 62176 25740 62240
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62176 26322 62240
rect 25702 62160 26322 62176
rect 25702 62096 25740 62160
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62096 26322 62160
rect 25702 62080 26322 62096
rect 25702 62016 25740 62080
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62016 26322 62080
rect 25702 62000 26322 62016
rect 25702 61936 25740 62000
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61936 26322 62000
rect 25702 52240 26322 61936
rect 25702 52176 25740 52240
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52176 26322 52240
rect 25702 52160 26322 52176
rect 25702 52096 25740 52160
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52096 26322 52160
rect 25702 52080 26322 52096
rect 25702 52016 25740 52080
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52016 26322 52080
rect 25702 52000 26322 52016
rect 25702 51936 25740 52000
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51936 26322 52000
rect 25702 42240 26322 51936
rect 25702 42176 25740 42240
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42176 26322 42240
rect 25702 42160 26322 42176
rect 25702 42096 25740 42160
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42096 26322 42160
rect 25702 42080 26322 42096
rect 25702 42016 25740 42080
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42016 26322 42080
rect 25702 42000 26322 42016
rect 25702 41936 25740 42000
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41936 26322 42000
rect 25702 32240 26322 41936
rect 25702 32176 25740 32240
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32176 26322 32240
rect 25702 32160 26322 32176
rect 25702 32096 25740 32160
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32096 26322 32160
rect 25702 32080 26322 32096
rect 25702 32016 25740 32080
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32016 26322 32080
rect 25702 32000 26322 32016
rect 25702 31936 25740 32000
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31936 26322 32000
rect 25702 22240 26322 31936
rect 25702 22176 25740 22240
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22176 26322 22240
rect 25702 22160 26322 22176
rect 25702 22096 25740 22160
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22096 26322 22160
rect 25702 22080 26322 22096
rect 25702 22016 25740 22080
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22016 26322 22080
rect 25702 22000 26322 22016
rect 25702 21936 25740 22000
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21936 26322 22000
rect 25702 12240 26322 21936
rect 25702 12176 25740 12240
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12176 26322 12240
rect 25702 12160 26322 12176
rect 25702 12096 25740 12160
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12096 26322 12160
rect 25702 12080 26322 12096
rect 25702 12016 25740 12080
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12016 26322 12080
rect 25702 12000 26322 12016
rect 25702 11936 25740 12000
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11936 26322 12000
rect 25702 2240 26322 11936
rect 25702 2176 25740 2240
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 26322 2240
rect 25702 2160 26322 2176
rect 25702 2096 25740 2160
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 26322 2160
rect 25702 2080 26322 2096
rect 25702 2016 25740 2080
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 26322 2080
rect 25702 2000 26322 2016
rect 25702 1936 25740 2000
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 26322 2000
rect 25702 0 26322 1936
rect 28702 84592 29322 87000
rect 28702 84528 28740 84592
rect 28804 84528 28820 84592
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84528 29322 84592
rect 28702 84512 29322 84528
rect 28702 84448 28740 84512
rect 28804 84448 28820 84512
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84448 29322 84512
rect 28702 84432 29322 84448
rect 28702 84368 28740 84432
rect 28804 84368 28820 84432
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84368 29322 84432
rect 28702 84352 29322 84368
rect 28702 84288 28740 84352
rect 28804 84288 28820 84352
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84288 29322 84352
rect 28702 74592 29322 84288
rect 28702 74528 28740 74592
rect 28804 74528 28820 74592
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74528 29322 74592
rect 28702 74512 29322 74528
rect 28702 74448 28740 74512
rect 28804 74448 28820 74512
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74448 29322 74512
rect 28702 74432 29322 74448
rect 28702 74368 28740 74432
rect 28804 74368 28820 74432
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74368 29322 74432
rect 28702 74352 29322 74368
rect 28702 74288 28740 74352
rect 28804 74288 28820 74352
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74288 29322 74352
rect 28702 64592 29322 74288
rect 28702 64528 28740 64592
rect 28804 64528 28820 64592
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64528 29322 64592
rect 28702 64512 29322 64528
rect 28702 64448 28740 64512
rect 28804 64448 28820 64512
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64448 29322 64512
rect 28702 64432 29322 64448
rect 28702 64368 28740 64432
rect 28804 64368 28820 64432
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64368 29322 64432
rect 28702 64352 29322 64368
rect 28702 64288 28740 64352
rect 28804 64288 28820 64352
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64288 29322 64352
rect 28702 54592 29322 64288
rect 28702 54528 28740 54592
rect 28804 54528 28820 54592
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54528 29322 54592
rect 28702 54512 29322 54528
rect 28702 54448 28740 54512
rect 28804 54448 28820 54512
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54448 29322 54512
rect 28702 54432 29322 54448
rect 28702 54368 28740 54432
rect 28804 54368 28820 54432
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54368 29322 54432
rect 28702 54352 29322 54368
rect 28702 54288 28740 54352
rect 28804 54288 28820 54352
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54288 29322 54352
rect 28702 44592 29322 54288
rect 28702 44528 28740 44592
rect 28804 44528 28820 44592
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44528 29322 44592
rect 28702 44512 29322 44528
rect 28702 44448 28740 44512
rect 28804 44448 28820 44512
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44448 29322 44512
rect 28702 44432 29322 44448
rect 28702 44368 28740 44432
rect 28804 44368 28820 44432
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44368 29322 44432
rect 28702 44352 29322 44368
rect 28702 44288 28740 44352
rect 28804 44288 28820 44352
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44288 29322 44352
rect 28702 34592 29322 44288
rect 28702 34528 28740 34592
rect 28804 34528 28820 34592
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34528 29322 34592
rect 28702 34512 29322 34528
rect 28702 34448 28740 34512
rect 28804 34448 28820 34512
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34448 29322 34512
rect 28702 34432 29322 34448
rect 28702 34368 28740 34432
rect 28804 34368 28820 34432
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34368 29322 34432
rect 28702 34352 29322 34368
rect 28702 34288 28740 34352
rect 28804 34288 28820 34352
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34288 29322 34352
rect 28702 24592 29322 34288
rect 28702 24528 28740 24592
rect 28804 24528 28820 24592
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24528 29322 24592
rect 28702 24512 29322 24528
rect 28702 24448 28740 24512
rect 28804 24448 28820 24512
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24448 29322 24512
rect 28702 24432 29322 24448
rect 28702 24368 28740 24432
rect 28804 24368 28820 24432
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24368 29322 24432
rect 28702 24352 29322 24368
rect 28702 24288 28740 24352
rect 28804 24288 28820 24352
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24288 29322 24352
rect 28702 14592 29322 24288
rect 28702 14528 28740 14592
rect 28804 14528 28820 14592
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14528 29322 14592
rect 28702 14512 29322 14528
rect 28702 14448 28740 14512
rect 28804 14448 28820 14512
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14448 29322 14512
rect 28702 14432 29322 14448
rect 28702 14368 28740 14432
rect 28804 14368 28820 14432
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14368 29322 14432
rect 28702 14352 29322 14368
rect 28702 14288 28740 14352
rect 28804 14288 28820 14352
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14288 29322 14352
rect 28702 4592 29322 14288
rect 28702 4528 28740 4592
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4528 29322 4592
rect 28702 4512 29322 4528
rect 28702 4448 28740 4512
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4448 29322 4512
rect 28702 4432 29322 4448
rect 28702 4368 28740 4432
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4368 29322 4432
rect 28702 4352 29322 4368
rect 28702 4288 28740 4352
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4288 29322 4352
rect 28702 0 29322 4288
rect 31702 82240 32322 87000
rect 31702 82176 31740 82240
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82176 32322 82240
rect 31702 82160 32322 82176
rect 31702 82096 31740 82160
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82096 32322 82160
rect 31702 82080 32322 82096
rect 31702 82016 31740 82080
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82016 32322 82080
rect 31702 82000 32322 82016
rect 31702 81936 31740 82000
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81936 32322 82000
rect 31702 72240 32322 81936
rect 31702 72176 31740 72240
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72176 32322 72240
rect 31702 72160 32322 72176
rect 31702 72096 31740 72160
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72096 32322 72160
rect 31702 72080 32322 72096
rect 31702 72016 31740 72080
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72016 32322 72080
rect 31702 72000 32322 72016
rect 31702 71936 31740 72000
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71936 32322 72000
rect 31702 62240 32322 71936
rect 31702 62176 31740 62240
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62176 32322 62240
rect 31702 62160 32322 62176
rect 31702 62096 31740 62160
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62096 32322 62160
rect 31702 62080 32322 62096
rect 31702 62016 31740 62080
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62016 32322 62080
rect 31702 62000 32322 62016
rect 31702 61936 31740 62000
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61936 32322 62000
rect 31702 52240 32322 61936
rect 31702 52176 31740 52240
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52176 32322 52240
rect 31702 52160 32322 52176
rect 31702 52096 31740 52160
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52096 32322 52160
rect 31702 52080 32322 52096
rect 31702 52016 31740 52080
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52016 32322 52080
rect 31702 52000 32322 52016
rect 31702 51936 31740 52000
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51936 32322 52000
rect 31702 42240 32322 51936
rect 31702 42176 31740 42240
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42176 32322 42240
rect 31702 42160 32322 42176
rect 31702 42096 31740 42160
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42096 32322 42160
rect 31702 42080 32322 42096
rect 31702 42016 31740 42080
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42016 32322 42080
rect 31702 42000 32322 42016
rect 31702 41936 31740 42000
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41936 32322 42000
rect 31702 32240 32322 41936
rect 31702 32176 31740 32240
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32176 32322 32240
rect 31702 32160 32322 32176
rect 31702 32096 31740 32160
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32096 32322 32160
rect 31702 32080 32322 32096
rect 31702 32016 31740 32080
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32016 32322 32080
rect 31702 32000 32322 32016
rect 31702 31936 31740 32000
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31936 32322 32000
rect 31702 22240 32322 31936
rect 31702 22176 31740 22240
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22176 32322 22240
rect 31702 22160 32322 22176
rect 31702 22096 31740 22160
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22096 32322 22160
rect 31702 22080 32322 22096
rect 31702 22016 31740 22080
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22016 32322 22080
rect 31702 22000 32322 22016
rect 31702 21936 31740 22000
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21936 32322 22000
rect 31702 12240 32322 21936
rect 31702 12176 31740 12240
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12176 32322 12240
rect 31702 12160 32322 12176
rect 31702 12096 31740 12160
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12096 32322 12160
rect 31702 12080 32322 12096
rect 31702 12016 31740 12080
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12016 32322 12080
rect 31702 12000 32322 12016
rect 31702 11936 31740 12000
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 32322 12000
rect 31702 2240 32322 11936
rect 31702 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2176 31900 2240
rect 31964 2176 31980 2240
rect 32044 2176 32060 2240
rect 32124 2176 32140 2240
rect 32204 2176 32220 2240
rect 32284 2176 32322 2240
rect 31702 2160 32322 2176
rect 31702 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2096 31900 2160
rect 31964 2096 31980 2160
rect 32044 2096 32060 2160
rect 32124 2096 32140 2160
rect 32204 2096 32220 2160
rect 32284 2096 32322 2160
rect 31702 2080 32322 2096
rect 31702 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2016 31900 2080
rect 31964 2016 31980 2080
rect 32044 2016 32060 2080
rect 32124 2016 32140 2080
rect 32204 2016 32220 2080
rect 32284 2016 32322 2080
rect 31702 2000 32322 2016
rect 31702 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1936 31900 2000
rect 31964 1936 31980 2000
rect 32044 1936 32060 2000
rect 32124 1936 32140 2000
rect 32204 1936 32220 2000
rect 32284 1936 32322 2000
rect 31702 0 32322 1936
rect 34702 84592 35322 87000
rect 34702 84528 34740 84592
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84528 35322 84592
rect 34702 84512 35322 84528
rect 34702 84448 34740 84512
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84448 35322 84512
rect 34702 84432 35322 84448
rect 34702 84368 34740 84432
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84368 35322 84432
rect 34702 84352 35322 84368
rect 34702 84288 34740 84352
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84288 35322 84352
rect 34702 74592 35322 84288
rect 34702 74528 34740 74592
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74528 35322 74592
rect 34702 74512 35322 74528
rect 34702 74448 34740 74512
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74448 35322 74512
rect 34702 74432 35322 74448
rect 34702 74368 34740 74432
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74368 35322 74432
rect 34702 74352 35322 74368
rect 34702 74288 34740 74352
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74288 35322 74352
rect 34702 64592 35322 74288
rect 34702 64528 34740 64592
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64528 35322 64592
rect 34702 64512 35322 64528
rect 34702 64448 34740 64512
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64448 35322 64512
rect 34702 64432 35322 64448
rect 34702 64368 34740 64432
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64368 35322 64432
rect 34702 64352 35322 64368
rect 34702 64288 34740 64352
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64288 35322 64352
rect 34702 54592 35322 64288
rect 34702 54528 34740 54592
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54528 35322 54592
rect 34702 54512 35322 54528
rect 34702 54448 34740 54512
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54448 35322 54512
rect 34702 54432 35322 54448
rect 34702 54368 34740 54432
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54368 35322 54432
rect 34702 54352 35322 54368
rect 34702 54288 34740 54352
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54288 35322 54352
rect 34702 44592 35322 54288
rect 34702 44528 34740 44592
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44528 35322 44592
rect 34702 44512 35322 44528
rect 34702 44448 34740 44512
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44448 35322 44512
rect 34702 44432 35322 44448
rect 34702 44368 34740 44432
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44368 35322 44432
rect 34702 44352 35322 44368
rect 34702 44288 34740 44352
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44288 35322 44352
rect 34702 34592 35322 44288
rect 34702 34528 34740 34592
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34528 35322 34592
rect 34702 34512 35322 34528
rect 34702 34448 34740 34512
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34448 35322 34512
rect 34702 34432 35322 34448
rect 34702 34368 34740 34432
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34368 35322 34432
rect 34702 34352 35322 34368
rect 34702 34288 34740 34352
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34288 35322 34352
rect 34702 24592 35322 34288
rect 34702 24528 34740 24592
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24528 35322 24592
rect 34702 24512 35322 24528
rect 34702 24448 34740 24512
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24448 35322 24512
rect 34702 24432 35322 24448
rect 34702 24368 34740 24432
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24368 35322 24432
rect 34702 24352 35322 24368
rect 34702 24288 34740 24352
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24288 35322 24352
rect 34702 14592 35322 24288
rect 34702 14528 34740 14592
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14528 35322 14592
rect 34702 14512 35322 14528
rect 34702 14448 34740 14512
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14448 35322 14512
rect 34702 14432 35322 14448
rect 34702 14368 34740 14432
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14368 35322 14432
rect 34702 14352 35322 14368
rect 34702 14288 34740 14352
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14288 35322 14352
rect 34702 4592 35322 14288
rect 34702 4528 34740 4592
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 35322 4592
rect 34702 4512 35322 4528
rect 34702 4448 34740 4512
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 35322 4512
rect 34702 4432 35322 4448
rect 34702 4368 34740 4432
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 35322 4432
rect 34702 4352 35322 4368
rect 34702 4288 34740 4352
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 35322 4352
rect 34702 0 35322 4288
rect 37702 82240 38322 87000
rect 37702 82176 37740 82240
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82176 38322 82240
rect 37702 82160 38322 82176
rect 37702 82096 37740 82160
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82096 38322 82160
rect 37702 82080 38322 82096
rect 37702 82016 37740 82080
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82016 38322 82080
rect 37702 82000 38322 82016
rect 37702 81936 37740 82000
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81936 38322 82000
rect 37702 72240 38322 81936
rect 37702 72176 37740 72240
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72176 38322 72240
rect 37702 72160 38322 72176
rect 37702 72096 37740 72160
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72096 38322 72160
rect 37702 72080 38322 72096
rect 37702 72016 37740 72080
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72016 38322 72080
rect 37702 72000 38322 72016
rect 37702 71936 37740 72000
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71936 38322 72000
rect 37702 62240 38322 71936
rect 37702 62176 37740 62240
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62176 38322 62240
rect 37702 62160 38322 62176
rect 37702 62096 37740 62160
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62096 38322 62160
rect 37702 62080 38322 62096
rect 37702 62016 37740 62080
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62016 38322 62080
rect 37702 62000 38322 62016
rect 37702 61936 37740 62000
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61936 38322 62000
rect 37702 52240 38322 61936
rect 37702 52176 37740 52240
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52176 38322 52240
rect 37702 52160 38322 52176
rect 37702 52096 37740 52160
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52096 38322 52160
rect 37702 52080 38322 52096
rect 37702 52016 37740 52080
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52016 38322 52080
rect 37702 52000 38322 52016
rect 37702 51936 37740 52000
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51936 38322 52000
rect 37702 42240 38322 51936
rect 37702 42176 37740 42240
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42176 38322 42240
rect 37702 42160 38322 42176
rect 37702 42096 37740 42160
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42096 38322 42160
rect 37702 42080 38322 42096
rect 37702 42016 37740 42080
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42016 38322 42080
rect 37702 42000 38322 42016
rect 37702 41936 37740 42000
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41936 38322 42000
rect 37702 32240 38322 41936
rect 37702 32176 37740 32240
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32176 38322 32240
rect 37702 32160 38322 32176
rect 37702 32096 37740 32160
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32096 38322 32160
rect 37702 32080 38322 32096
rect 37702 32016 37740 32080
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32016 38322 32080
rect 37702 32000 38322 32016
rect 37702 31936 37740 32000
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31936 38322 32000
rect 37702 22240 38322 31936
rect 37702 22176 37740 22240
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22176 38322 22240
rect 37702 22160 38322 22176
rect 37702 22096 37740 22160
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22096 38322 22160
rect 37702 22080 38322 22096
rect 37702 22016 37740 22080
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22016 38322 22080
rect 37702 22000 38322 22016
rect 37702 21936 37740 22000
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21936 38322 22000
rect 37702 12240 38322 21936
rect 37702 12176 37740 12240
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12176 38322 12240
rect 37702 12160 38322 12176
rect 37702 12096 37740 12160
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12096 38322 12160
rect 37702 12080 38322 12096
rect 37702 12016 37740 12080
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12016 38322 12080
rect 37702 12000 38322 12016
rect 37702 11936 37740 12000
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11936 38322 12000
rect 37702 2240 38322 11936
rect 40702 84592 41322 87000
rect 40702 84528 40740 84592
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84528 41322 84592
rect 40702 84512 41322 84528
rect 40702 84448 40740 84512
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84448 41322 84512
rect 40702 84432 41322 84448
rect 40702 84368 40740 84432
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84368 41322 84432
rect 40702 84352 41322 84368
rect 40702 84288 40740 84352
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84288 41322 84352
rect 40702 74592 41322 84288
rect 40702 74528 40740 74592
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74528 41322 74592
rect 40702 74512 41322 74528
rect 40702 74448 40740 74512
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74448 41322 74512
rect 40702 74432 41322 74448
rect 40702 74368 40740 74432
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74368 41322 74432
rect 40702 74352 41322 74368
rect 40702 74288 40740 74352
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74288 41322 74352
rect 40702 64592 41322 74288
rect 40702 64528 40740 64592
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64528 41322 64592
rect 40702 64512 41322 64528
rect 40702 64448 40740 64512
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64448 41322 64512
rect 40702 64432 41322 64448
rect 40702 64368 40740 64432
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64368 41322 64432
rect 40702 64352 41322 64368
rect 40702 64288 40740 64352
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64288 41322 64352
rect 40702 54592 41322 64288
rect 40702 54528 40740 54592
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54528 41322 54592
rect 40702 54512 41322 54528
rect 40702 54448 40740 54512
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54448 41322 54512
rect 40702 54432 41322 54448
rect 40702 54368 40740 54432
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54368 41322 54432
rect 40702 54352 41322 54368
rect 40702 54288 40740 54352
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54288 41322 54352
rect 40702 44592 41322 54288
rect 40702 44528 40740 44592
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44528 41322 44592
rect 40702 44512 41322 44528
rect 40702 44448 40740 44512
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44448 41322 44512
rect 40702 44432 41322 44448
rect 40702 44368 40740 44432
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44368 41322 44432
rect 40702 44352 41322 44368
rect 40702 44288 40740 44352
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44288 41322 44352
rect 40702 34592 41322 44288
rect 40702 34528 40740 34592
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34528 41322 34592
rect 40702 34512 41322 34528
rect 40702 34448 40740 34512
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34448 41322 34512
rect 40702 34432 41322 34448
rect 40702 34368 40740 34432
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34368 41322 34432
rect 40702 34352 41322 34368
rect 40702 34288 40740 34352
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34288 41322 34352
rect 40702 24592 41322 34288
rect 40702 24528 40740 24592
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24528 41322 24592
rect 40702 24512 41322 24528
rect 40702 24448 40740 24512
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24448 41322 24512
rect 40702 24432 41322 24448
rect 40702 24368 40740 24432
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24368 41322 24432
rect 40702 24352 41322 24368
rect 40702 24288 40740 24352
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24288 41322 24352
rect 40702 14592 41322 24288
rect 40702 14528 40740 14592
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14528 41322 14592
rect 40702 14512 41322 14528
rect 40702 14448 40740 14512
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14448 41322 14512
rect 40702 14432 41322 14448
rect 40702 14368 40740 14432
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14368 41322 14432
rect 40702 14352 41322 14368
rect 40702 14288 40740 14352
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14288 41322 14352
rect 39987 5812 40053 5813
rect 39987 5748 39988 5812
rect 40052 5748 40053 5812
rect 39987 5747 40053 5748
rect 39990 3365 40050 5747
rect 40702 4592 41322 14288
rect 40702 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4528 41322 4592
rect 40702 4512 41322 4528
rect 40702 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4448 41322 4512
rect 40702 4432 41322 4448
rect 40702 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4368 41322 4432
rect 40702 4352 41322 4368
rect 40702 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4288 41322 4352
rect 39987 3364 40053 3365
rect 39987 3300 39988 3364
rect 40052 3300 40053 3364
rect 39987 3299 40053 3300
rect 37702 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2176 38322 2240
rect 37702 2160 38322 2176
rect 37702 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2096 38322 2160
rect 37702 2080 38322 2096
rect 37702 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2016 38322 2080
rect 37702 2000 38322 2016
rect 37702 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1936 38322 2000
rect 37702 0 38322 1936
rect 40702 0 41322 4288
rect 43702 82240 44322 87000
rect 43702 82176 43740 82240
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82176 44322 82240
rect 43702 82160 44322 82176
rect 43702 82096 43740 82160
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82096 44322 82160
rect 43702 82080 44322 82096
rect 43702 82016 43740 82080
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82016 44322 82080
rect 43702 82000 44322 82016
rect 43702 81936 43740 82000
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81936 44322 82000
rect 43702 72240 44322 81936
rect 43702 72176 43740 72240
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72176 44322 72240
rect 43702 72160 44322 72176
rect 43702 72096 43740 72160
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72096 44322 72160
rect 43702 72080 44322 72096
rect 43702 72016 43740 72080
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72016 44322 72080
rect 43702 72000 44322 72016
rect 43702 71936 43740 72000
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71936 44322 72000
rect 43702 62240 44322 71936
rect 43702 62176 43740 62240
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62176 44322 62240
rect 43702 62160 44322 62176
rect 43702 62096 43740 62160
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62096 44322 62160
rect 43702 62080 44322 62096
rect 43702 62016 43740 62080
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62016 44322 62080
rect 43702 62000 44322 62016
rect 43702 61936 43740 62000
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61936 44322 62000
rect 43702 52240 44322 61936
rect 43702 52176 43740 52240
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52176 44322 52240
rect 43702 52160 44322 52176
rect 43702 52096 43740 52160
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52096 44322 52160
rect 43702 52080 44322 52096
rect 43702 52016 43740 52080
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52016 44322 52080
rect 43702 52000 44322 52016
rect 43702 51936 43740 52000
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51936 44322 52000
rect 43702 42240 44322 51936
rect 43702 42176 43740 42240
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42176 44322 42240
rect 43702 42160 44322 42176
rect 43702 42096 43740 42160
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42096 44322 42160
rect 43702 42080 44322 42096
rect 43702 42016 43740 42080
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42016 44322 42080
rect 43702 42000 44322 42016
rect 43702 41936 43740 42000
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41936 44322 42000
rect 43702 32240 44322 41936
rect 43702 32176 43740 32240
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32176 44322 32240
rect 43702 32160 44322 32176
rect 43702 32096 43740 32160
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32096 44322 32160
rect 43702 32080 44322 32096
rect 43702 32016 43740 32080
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32016 44322 32080
rect 43702 32000 44322 32016
rect 43702 31936 43740 32000
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31936 44322 32000
rect 43702 22240 44322 31936
rect 43702 22176 43740 22240
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22176 44322 22240
rect 43702 22160 44322 22176
rect 43702 22096 43740 22160
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22096 44322 22160
rect 43702 22080 44322 22096
rect 43702 22016 43740 22080
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22016 44322 22080
rect 43702 22000 44322 22016
rect 43702 21936 43740 22000
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21936 44322 22000
rect 43702 12240 44322 21936
rect 43702 12176 43740 12240
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12176 44322 12240
rect 43702 12160 44322 12176
rect 43702 12096 43740 12160
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12096 44322 12160
rect 43702 12080 44322 12096
rect 43702 12016 43740 12080
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12016 44322 12080
rect 43702 12000 44322 12016
rect 43702 11936 43740 12000
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11936 44322 12000
rect 43702 2240 44322 11936
rect 43702 2176 43740 2240
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 44322 2240
rect 43702 2160 44322 2176
rect 43702 2096 43740 2160
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 44322 2160
rect 43702 2080 44322 2096
rect 43702 2016 43740 2080
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 44322 2080
rect 43702 2000 44322 2016
rect 43702 1936 43740 2000
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 44322 2000
rect 43702 0 44322 1936
rect 46702 84592 47322 87000
rect 46702 84528 46740 84592
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84528 47322 84592
rect 46702 84512 47322 84528
rect 46702 84448 46740 84512
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84448 47322 84512
rect 46702 84432 47322 84448
rect 46702 84368 46740 84432
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84368 47322 84432
rect 46702 84352 47322 84368
rect 46702 84288 46740 84352
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84288 47322 84352
rect 46702 74592 47322 84288
rect 46702 74528 46740 74592
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74528 47322 74592
rect 46702 74512 47322 74528
rect 46702 74448 46740 74512
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74448 47322 74512
rect 46702 74432 47322 74448
rect 46702 74368 46740 74432
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74368 47322 74432
rect 46702 74352 47322 74368
rect 46702 74288 46740 74352
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74288 47322 74352
rect 46702 64592 47322 74288
rect 46702 64528 46740 64592
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64528 47322 64592
rect 46702 64512 47322 64528
rect 46702 64448 46740 64512
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64448 47322 64512
rect 46702 64432 47322 64448
rect 46702 64368 46740 64432
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64368 47322 64432
rect 46702 64352 47322 64368
rect 46702 64288 46740 64352
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64288 47322 64352
rect 46702 54592 47322 64288
rect 46702 54528 46740 54592
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54528 47322 54592
rect 46702 54512 47322 54528
rect 46702 54448 46740 54512
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54448 47322 54512
rect 46702 54432 47322 54448
rect 46702 54368 46740 54432
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54368 47322 54432
rect 46702 54352 47322 54368
rect 46702 54288 46740 54352
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54288 47322 54352
rect 46702 44592 47322 54288
rect 46702 44528 46740 44592
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44528 47322 44592
rect 46702 44512 47322 44528
rect 46702 44448 46740 44512
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44448 47322 44512
rect 46702 44432 47322 44448
rect 46702 44368 46740 44432
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44368 47322 44432
rect 46702 44352 47322 44368
rect 46702 44288 46740 44352
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44288 47322 44352
rect 46702 34592 47322 44288
rect 46702 34528 46740 34592
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34528 47322 34592
rect 46702 34512 47322 34528
rect 46702 34448 46740 34512
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34448 47322 34512
rect 46702 34432 47322 34448
rect 46702 34368 46740 34432
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34368 47322 34432
rect 46702 34352 47322 34368
rect 46702 34288 46740 34352
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34288 47322 34352
rect 46702 24592 47322 34288
rect 46702 24528 46740 24592
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24528 47322 24592
rect 46702 24512 47322 24528
rect 46702 24448 46740 24512
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24448 47322 24512
rect 46702 24432 47322 24448
rect 46702 24368 46740 24432
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24368 47322 24432
rect 46702 24352 47322 24368
rect 46702 24288 46740 24352
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24288 47322 24352
rect 46702 14592 47322 24288
rect 46702 14528 46740 14592
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14528 47322 14592
rect 46702 14512 47322 14528
rect 46702 14448 46740 14512
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14448 47322 14512
rect 46702 14432 47322 14448
rect 46702 14368 46740 14432
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14368 47322 14432
rect 46702 14352 47322 14368
rect 46702 14288 46740 14352
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14288 47322 14352
rect 46702 4592 47322 14288
rect 46702 4528 46740 4592
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 47322 4592
rect 46702 4512 47322 4528
rect 46702 4448 46740 4512
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 47322 4512
rect 46702 4432 47322 4448
rect 46702 4368 46740 4432
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 47322 4432
rect 46702 4352 47322 4368
rect 46702 4288 46740 4352
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 47322 4352
rect 46702 0 47322 4288
rect 49702 82240 50322 87000
rect 49702 82176 49740 82240
rect 49804 82176 49820 82240
rect 49884 82176 49900 82240
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82176 50322 82240
rect 49702 82160 50322 82176
rect 49702 82096 49740 82160
rect 49804 82096 49820 82160
rect 49884 82096 49900 82160
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82096 50322 82160
rect 49702 82080 50322 82096
rect 49702 82016 49740 82080
rect 49804 82016 49820 82080
rect 49884 82016 49900 82080
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82016 50322 82080
rect 49702 82000 50322 82016
rect 49702 81936 49740 82000
rect 49804 81936 49820 82000
rect 49884 81936 49900 82000
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81936 50322 82000
rect 49702 72240 50322 81936
rect 49702 72176 49740 72240
rect 49804 72176 49820 72240
rect 49884 72176 49900 72240
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72176 50322 72240
rect 49702 72160 50322 72176
rect 49702 72096 49740 72160
rect 49804 72096 49820 72160
rect 49884 72096 49900 72160
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72096 50322 72160
rect 49702 72080 50322 72096
rect 49702 72016 49740 72080
rect 49804 72016 49820 72080
rect 49884 72016 49900 72080
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72016 50322 72080
rect 49702 72000 50322 72016
rect 49702 71936 49740 72000
rect 49804 71936 49820 72000
rect 49884 71936 49900 72000
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71936 50322 72000
rect 49702 62240 50322 71936
rect 49702 62176 49740 62240
rect 49804 62176 49820 62240
rect 49884 62176 49900 62240
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62176 50322 62240
rect 49702 62160 50322 62176
rect 49702 62096 49740 62160
rect 49804 62096 49820 62160
rect 49884 62096 49900 62160
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62096 50322 62160
rect 49702 62080 50322 62096
rect 49702 62016 49740 62080
rect 49804 62016 49820 62080
rect 49884 62016 49900 62080
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62016 50322 62080
rect 49702 62000 50322 62016
rect 49702 61936 49740 62000
rect 49804 61936 49820 62000
rect 49884 61936 49900 62000
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61936 50322 62000
rect 49702 52240 50322 61936
rect 49702 52176 49740 52240
rect 49804 52176 49820 52240
rect 49884 52176 49900 52240
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52176 50322 52240
rect 49702 52160 50322 52176
rect 49702 52096 49740 52160
rect 49804 52096 49820 52160
rect 49884 52096 49900 52160
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52096 50322 52160
rect 49702 52080 50322 52096
rect 49702 52016 49740 52080
rect 49804 52016 49820 52080
rect 49884 52016 49900 52080
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52016 50322 52080
rect 49702 52000 50322 52016
rect 49702 51936 49740 52000
rect 49804 51936 49820 52000
rect 49884 51936 49900 52000
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51936 50322 52000
rect 49702 42240 50322 51936
rect 49702 42176 49740 42240
rect 49804 42176 49820 42240
rect 49884 42176 49900 42240
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42176 50322 42240
rect 49702 42160 50322 42176
rect 49702 42096 49740 42160
rect 49804 42096 49820 42160
rect 49884 42096 49900 42160
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42096 50322 42160
rect 49702 42080 50322 42096
rect 49702 42016 49740 42080
rect 49804 42016 49820 42080
rect 49884 42016 49900 42080
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42016 50322 42080
rect 49702 42000 50322 42016
rect 49702 41936 49740 42000
rect 49804 41936 49820 42000
rect 49884 41936 49900 42000
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41936 50322 42000
rect 49702 32240 50322 41936
rect 49702 32176 49740 32240
rect 49804 32176 49820 32240
rect 49884 32176 49900 32240
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32176 50322 32240
rect 49702 32160 50322 32176
rect 49702 32096 49740 32160
rect 49804 32096 49820 32160
rect 49884 32096 49900 32160
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32096 50322 32160
rect 49702 32080 50322 32096
rect 49702 32016 49740 32080
rect 49804 32016 49820 32080
rect 49884 32016 49900 32080
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32016 50322 32080
rect 49702 32000 50322 32016
rect 49702 31936 49740 32000
rect 49804 31936 49820 32000
rect 49884 31936 49900 32000
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31936 50322 32000
rect 49702 22240 50322 31936
rect 49702 22176 49740 22240
rect 49804 22176 49820 22240
rect 49884 22176 49900 22240
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22176 50322 22240
rect 49702 22160 50322 22176
rect 49702 22096 49740 22160
rect 49804 22096 49820 22160
rect 49884 22096 49900 22160
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22096 50322 22160
rect 49702 22080 50322 22096
rect 49702 22016 49740 22080
rect 49804 22016 49820 22080
rect 49884 22016 49900 22080
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22016 50322 22080
rect 49702 22000 50322 22016
rect 49702 21936 49740 22000
rect 49804 21936 49820 22000
rect 49884 21936 49900 22000
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21936 50322 22000
rect 49702 12240 50322 21936
rect 49702 12176 49740 12240
rect 49804 12176 49820 12240
rect 49884 12176 49900 12240
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12176 50322 12240
rect 49702 12160 50322 12176
rect 49702 12096 49740 12160
rect 49804 12096 49820 12160
rect 49884 12096 49900 12160
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12096 50322 12160
rect 49702 12080 50322 12096
rect 49702 12016 49740 12080
rect 49804 12016 49820 12080
rect 49884 12016 49900 12080
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12016 50322 12080
rect 49702 12000 50322 12016
rect 49702 11936 49740 12000
rect 49804 11936 49820 12000
rect 49884 11936 49900 12000
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11936 50322 12000
rect 49702 2240 50322 11936
rect 49702 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2176 50322 2240
rect 49702 2160 50322 2176
rect 49702 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2096 50322 2160
rect 49702 2080 50322 2096
rect 49702 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2016 50322 2080
rect 49702 2000 50322 2016
rect 49702 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1936 50322 2000
rect 49702 0 50322 1936
rect 52702 84592 53322 87000
rect 52702 84528 52740 84592
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84528 53322 84592
rect 52702 84512 53322 84528
rect 52702 84448 52740 84512
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84448 53322 84512
rect 52702 84432 53322 84448
rect 52702 84368 52740 84432
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84368 53322 84432
rect 52702 84352 53322 84368
rect 52702 84288 52740 84352
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84288 53322 84352
rect 52702 74592 53322 84288
rect 52702 74528 52740 74592
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74528 53322 74592
rect 52702 74512 53322 74528
rect 52702 74448 52740 74512
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74448 53322 74512
rect 52702 74432 53322 74448
rect 52702 74368 52740 74432
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74368 53322 74432
rect 52702 74352 53322 74368
rect 52702 74288 52740 74352
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74288 53322 74352
rect 52702 64592 53322 74288
rect 52702 64528 52740 64592
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64528 53322 64592
rect 52702 64512 53322 64528
rect 52702 64448 52740 64512
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64448 53322 64512
rect 52702 64432 53322 64448
rect 52702 64368 52740 64432
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64368 53322 64432
rect 52702 64352 53322 64368
rect 52702 64288 52740 64352
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64288 53322 64352
rect 52702 54592 53322 64288
rect 52702 54528 52740 54592
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54528 53322 54592
rect 52702 54512 53322 54528
rect 52702 54448 52740 54512
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54448 53322 54512
rect 52702 54432 53322 54448
rect 52702 54368 52740 54432
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54368 53322 54432
rect 52702 54352 53322 54368
rect 52702 54288 52740 54352
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54288 53322 54352
rect 52702 44592 53322 54288
rect 52702 44528 52740 44592
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44528 53322 44592
rect 52702 44512 53322 44528
rect 52702 44448 52740 44512
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44448 53322 44512
rect 52702 44432 53322 44448
rect 52702 44368 52740 44432
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44368 53322 44432
rect 52702 44352 53322 44368
rect 52702 44288 52740 44352
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44288 53322 44352
rect 52702 34592 53322 44288
rect 52702 34528 52740 34592
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34528 53322 34592
rect 52702 34512 53322 34528
rect 52702 34448 52740 34512
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34448 53322 34512
rect 52702 34432 53322 34448
rect 52702 34368 52740 34432
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34368 53322 34432
rect 52702 34352 53322 34368
rect 52702 34288 52740 34352
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34288 53322 34352
rect 52702 24592 53322 34288
rect 52702 24528 52740 24592
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24528 53322 24592
rect 52702 24512 53322 24528
rect 52702 24448 52740 24512
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24448 53322 24512
rect 52702 24432 53322 24448
rect 52702 24368 52740 24432
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24368 53322 24432
rect 52702 24352 53322 24368
rect 52702 24288 52740 24352
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24288 53322 24352
rect 52702 14592 53322 24288
rect 52702 14528 52740 14592
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14528 53322 14592
rect 52702 14512 53322 14528
rect 52702 14448 52740 14512
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14448 53322 14512
rect 52702 14432 53322 14448
rect 52702 14368 52740 14432
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14368 53322 14432
rect 52702 14352 53322 14368
rect 52702 14288 52740 14352
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14288 53322 14352
rect 52702 4592 53322 14288
rect 52702 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4528 53322 4592
rect 52702 4512 53322 4528
rect 52702 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4448 53322 4512
rect 52702 4432 53322 4448
rect 52702 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4368 53322 4432
rect 52702 4352 53322 4368
rect 52702 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4288 53322 4352
rect 52702 0 53322 4288
rect 55702 82240 56322 87000
rect 55702 82176 55740 82240
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82176 56322 82240
rect 55702 82160 56322 82176
rect 55702 82096 55740 82160
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82096 56322 82160
rect 55702 82080 56322 82096
rect 55702 82016 55740 82080
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82016 56322 82080
rect 55702 82000 56322 82016
rect 55702 81936 55740 82000
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81936 56322 82000
rect 55702 72240 56322 81936
rect 55702 72176 55740 72240
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72176 56322 72240
rect 55702 72160 56322 72176
rect 55702 72096 55740 72160
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72096 56322 72160
rect 55702 72080 56322 72096
rect 55702 72016 55740 72080
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72016 56322 72080
rect 55702 72000 56322 72016
rect 55702 71936 55740 72000
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71936 56322 72000
rect 55702 62240 56322 71936
rect 55702 62176 55740 62240
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62176 56322 62240
rect 55702 62160 56322 62176
rect 55702 62096 55740 62160
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62096 56322 62160
rect 55702 62080 56322 62096
rect 55702 62016 55740 62080
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62016 56322 62080
rect 55702 62000 56322 62016
rect 55702 61936 55740 62000
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61936 56322 62000
rect 55702 52240 56322 61936
rect 55702 52176 55740 52240
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52176 56322 52240
rect 55702 52160 56322 52176
rect 55702 52096 55740 52160
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52096 56322 52160
rect 55702 52080 56322 52096
rect 55702 52016 55740 52080
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52016 56322 52080
rect 55702 52000 56322 52016
rect 55702 51936 55740 52000
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51936 56322 52000
rect 55702 42240 56322 51936
rect 55702 42176 55740 42240
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42176 56322 42240
rect 55702 42160 56322 42176
rect 55702 42096 55740 42160
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42096 56322 42160
rect 55702 42080 56322 42096
rect 55702 42016 55740 42080
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42016 56322 42080
rect 55702 42000 56322 42016
rect 55702 41936 55740 42000
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41936 56322 42000
rect 55702 32240 56322 41936
rect 55702 32176 55740 32240
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32176 56322 32240
rect 55702 32160 56322 32176
rect 55702 32096 55740 32160
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32096 56322 32160
rect 55702 32080 56322 32096
rect 55702 32016 55740 32080
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32016 56322 32080
rect 55702 32000 56322 32016
rect 55702 31936 55740 32000
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31936 56322 32000
rect 55702 22240 56322 31936
rect 55702 22176 55740 22240
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22176 56322 22240
rect 55702 22160 56322 22176
rect 55702 22096 55740 22160
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22096 56322 22160
rect 55702 22080 56322 22096
rect 55702 22016 55740 22080
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22016 56322 22080
rect 55702 22000 56322 22016
rect 55702 21936 55740 22000
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21936 56322 22000
rect 55702 12240 56322 21936
rect 55702 12176 55740 12240
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12176 56322 12240
rect 55702 12160 56322 12176
rect 55702 12096 55740 12160
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12096 56322 12160
rect 55702 12080 56322 12096
rect 55702 12016 55740 12080
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12016 56322 12080
rect 55702 12000 56322 12016
rect 55702 11936 55740 12000
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11936 56322 12000
rect 55702 2240 56322 11936
rect 55702 2176 55740 2240
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 56322 2240
rect 55702 2160 56322 2176
rect 55702 2096 55740 2160
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 56322 2160
rect 55702 2080 56322 2096
rect 55702 2016 55740 2080
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 56322 2080
rect 55702 2000 56322 2016
rect 55702 1936 55740 2000
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 56322 2000
rect 55702 0 56322 1936
rect 58702 84592 59322 87000
rect 58702 84528 58740 84592
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84528 59060 84592
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84528 59322 84592
rect 58702 84512 59322 84528
rect 58702 84448 58740 84512
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84448 59060 84512
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84448 59322 84512
rect 58702 84432 59322 84448
rect 58702 84368 58740 84432
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84368 59060 84432
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84368 59322 84432
rect 58702 84352 59322 84368
rect 58702 84288 58740 84352
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84288 59060 84352
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84288 59322 84352
rect 58702 74592 59322 84288
rect 58702 74528 58740 74592
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74528 59060 74592
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74528 59322 74592
rect 58702 74512 59322 74528
rect 58702 74448 58740 74512
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74448 59060 74512
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74448 59322 74512
rect 58702 74432 59322 74448
rect 58702 74368 58740 74432
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74368 59060 74432
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74368 59322 74432
rect 58702 74352 59322 74368
rect 58702 74288 58740 74352
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74288 59060 74352
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74288 59322 74352
rect 58702 64592 59322 74288
rect 58702 64528 58740 64592
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64528 59060 64592
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64528 59322 64592
rect 58702 64512 59322 64528
rect 58702 64448 58740 64512
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64448 59060 64512
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64448 59322 64512
rect 58702 64432 59322 64448
rect 58702 64368 58740 64432
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64368 59060 64432
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64368 59322 64432
rect 58702 64352 59322 64368
rect 58702 64288 58740 64352
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64288 59060 64352
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64288 59322 64352
rect 58702 54592 59322 64288
rect 58702 54528 58740 54592
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54528 59060 54592
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54528 59322 54592
rect 58702 54512 59322 54528
rect 58702 54448 58740 54512
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54448 59060 54512
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54448 59322 54512
rect 58702 54432 59322 54448
rect 58702 54368 58740 54432
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54368 59060 54432
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54368 59322 54432
rect 58702 54352 59322 54368
rect 58702 54288 58740 54352
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54288 59060 54352
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54288 59322 54352
rect 58702 44592 59322 54288
rect 58702 44528 58740 44592
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44528 59060 44592
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44528 59322 44592
rect 58702 44512 59322 44528
rect 58702 44448 58740 44512
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44448 59060 44512
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44448 59322 44512
rect 58702 44432 59322 44448
rect 58702 44368 58740 44432
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44368 59060 44432
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44368 59322 44432
rect 58702 44352 59322 44368
rect 58702 44288 58740 44352
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44288 59060 44352
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44288 59322 44352
rect 58702 34592 59322 44288
rect 58702 34528 58740 34592
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34528 59060 34592
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34528 59322 34592
rect 58702 34512 59322 34528
rect 58702 34448 58740 34512
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34448 59060 34512
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34448 59322 34512
rect 58702 34432 59322 34448
rect 58702 34368 58740 34432
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34368 59060 34432
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34368 59322 34432
rect 58702 34352 59322 34368
rect 58702 34288 58740 34352
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34288 59060 34352
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34288 59322 34352
rect 58702 24592 59322 34288
rect 58702 24528 58740 24592
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24528 59060 24592
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24528 59322 24592
rect 58702 24512 59322 24528
rect 58702 24448 58740 24512
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24448 59060 24512
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24448 59322 24512
rect 58702 24432 59322 24448
rect 58702 24368 58740 24432
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24368 59060 24432
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24368 59322 24432
rect 58702 24352 59322 24368
rect 58702 24288 58740 24352
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24288 59060 24352
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24288 59322 24352
rect 58702 14592 59322 24288
rect 58702 14528 58740 14592
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14528 59060 14592
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14528 59322 14592
rect 58702 14512 59322 14528
rect 58702 14448 58740 14512
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14448 59060 14512
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14448 59322 14512
rect 58702 14432 59322 14448
rect 58702 14368 58740 14432
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14368 59060 14432
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14368 59322 14432
rect 58702 14352 59322 14368
rect 58702 14288 58740 14352
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14288 59060 14352
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14288 59322 14352
rect 58702 4592 59322 14288
rect 58702 4528 58740 4592
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4528 59322 4592
rect 58702 4512 59322 4528
rect 58702 4448 58740 4512
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4448 59322 4512
rect 58702 4432 59322 4448
rect 58702 4368 58740 4432
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4368 59322 4432
rect 58702 4352 59322 4368
rect 58702 4288 58740 4352
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4288 59322 4352
rect 58702 0 59322 4288
rect 61702 82240 62322 87000
rect 61702 82176 61740 82240
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82176 62322 82240
rect 61702 82160 62322 82176
rect 61702 82096 61740 82160
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82096 62322 82160
rect 61702 82080 62322 82096
rect 61702 82016 61740 82080
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82016 62322 82080
rect 61702 82000 62322 82016
rect 61702 81936 61740 82000
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81936 62322 82000
rect 61702 72240 62322 81936
rect 61702 72176 61740 72240
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72176 62322 72240
rect 61702 72160 62322 72176
rect 61702 72096 61740 72160
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72096 62322 72160
rect 61702 72080 62322 72096
rect 61702 72016 61740 72080
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72016 62322 72080
rect 61702 72000 62322 72016
rect 61702 71936 61740 72000
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71936 62322 72000
rect 61702 62240 62322 71936
rect 61702 62176 61740 62240
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62176 62322 62240
rect 61702 62160 62322 62176
rect 61702 62096 61740 62160
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62096 62322 62160
rect 61702 62080 62322 62096
rect 61702 62016 61740 62080
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62016 62322 62080
rect 61702 62000 62322 62016
rect 61702 61936 61740 62000
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61936 62322 62000
rect 61702 52240 62322 61936
rect 64702 84592 65322 87000
rect 64702 84528 64740 84592
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 65322 84592
rect 64702 84512 65322 84528
rect 64702 84448 64740 84512
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 65322 84512
rect 64702 84432 65322 84448
rect 64702 84368 64740 84432
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 65322 84432
rect 64702 84352 65322 84368
rect 64702 84288 64740 84352
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 65322 84352
rect 64702 74592 65322 84288
rect 64702 74528 64740 74592
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 65322 74592
rect 64702 74512 65322 74528
rect 64702 74448 64740 74512
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 65322 74512
rect 64702 74432 65322 74448
rect 64702 74368 64740 74432
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 65322 74432
rect 64702 74352 65322 74368
rect 64702 74288 64740 74352
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 65322 74352
rect 64702 64592 65322 74288
rect 64702 64528 64740 64592
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 65322 64592
rect 64702 64512 65322 64528
rect 64702 64448 64740 64512
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 65322 64512
rect 64702 64432 65322 64448
rect 64702 64368 64740 64432
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 65322 64432
rect 64702 64352 65322 64368
rect 64702 64288 64740 64352
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 65322 64352
rect 64702 54592 65322 64288
rect 64702 54528 64740 54592
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 65322 54592
rect 64702 54512 65322 54528
rect 64702 54448 64740 54512
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 65322 54512
rect 64702 54432 65322 54448
rect 64702 54368 64740 54432
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 65322 54432
rect 64702 54352 65322 54368
rect 64702 54288 64740 54352
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 65322 54352
rect 64091 52596 64157 52597
rect 64091 52532 64092 52596
rect 64156 52532 64157 52596
rect 64091 52531 64157 52532
rect 61702 52176 61740 52240
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52176 62322 52240
rect 61702 52160 62322 52176
rect 61702 52096 61740 52160
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52096 62322 52160
rect 61702 52080 62322 52096
rect 61702 52016 61740 52080
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52016 62322 52080
rect 61702 52000 62322 52016
rect 61702 51936 61740 52000
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51936 62322 52000
rect 61702 42240 62322 51936
rect 63171 44844 63237 44845
rect 63171 44780 63172 44844
rect 63236 44780 63237 44844
rect 63171 44779 63237 44780
rect 61702 42176 61740 42240
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42176 62322 42240
rect 61702 42160 62322 42176
rect 61702 42096 61740 42160
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42096 62322 42160
rect 61702 42080 62322 42096
rect 61702 42016 61740 42080
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42016 62322 42080
rect 61702 42000 62322 42016
rect 61702 41936 61740 42000
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41936 62322 42000
rect 61702 32240 62322 41936
rect 61702 32176 61740 32240
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32176 62322 32240
rect 61702 32160 62322 32176
rect 61702 32096 61740 32160
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32096 62322 32160
rect 61702 32080 62322 32096
rect 61702 32016 61740 32080
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32016 62322 32080
rect 61702 32000 62322 32016
rect 61702 31936 61740 32000
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31936 62322 32000
rect 61702 22240 62322 31936
rect 61702 22176 61740 22240
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22176 62322 22240
rect 61702 22160 62322 22176
rect 61702 22096 61740 22160
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22096 62322 22160
rect 61702 22080 62322 22096
rect 61702 22016 61740 22080
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22016 62322 22080
rect 61702 22000 62322 22016
rect 61702 21936 61740 22000
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21936 62322 22000
rect 61702 12240 62322 21936
rect 62987 17916 63053 17917
rect 62987 17852 62988 17916
rect 63052 17852 63053 17916
rect 62987 17851 63053 17852
rect 61702 12176 61740 12240
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12176 62322 12240
rect 61702 12160 62322 12176
rect 61702 12096 61740 12160
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12096 62322 12160
rect 61702 12080 62322 12096
rect 61702 12016 61740 12080
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12016 62322 12080
rect 61702 12000 62322 12016
rect 61702 11936 61740 12000
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11936 62322 12000
rect 61702 2240 62322 11936
rect 62990 6901 63050 17851
rect 62987 6900 63053 6901
rect 62987 6836 62988 6900
rect 63052 6836 63053 6900
rect 62987 6835 63053 6836
rect 63174 4861 63234 44779
rect 63907 43348 63973 43349
rect 63907 43284 63908 43348
rect 63972 43284 63973 43348
rect 63907 43283 63973 43284
rect 63723 12476 63789 12477
rect 63723 12412 63724 12476
rect 63788 12412 63789 12476
rect 63723 12411 63789 12412
rect 63726 11797 63786 12411
rect 63723 11796 63789 11797
rect 63723 11732 63724 11796
rect 63788 11732 63789 11796
rect 63723 11731 63789 11732
rect 63910 7717 63970 43283
rect 63907 7716 63973 7717
rect 63907 7652 63908 7716
rect 63972 7652 63973 7716
rect 63907 7651 63973 7652
rect 64094 5405 64154 52531
rect 64275 50284 64341 50285
rect 64275 50220 64276 50284
rect 64340 50220 64341 50284
rect 64275 50219 64341 50220
rect 64091 5404 64157 5405
rect 64091 5340 64092 5404
rect 64156 5340 64157 5404
rect 64091 5339 64157 5340
rect 64278 4997 64338 50219
rect 64459 47700 64525 47701
rect 64459 47636 64460 47700
rect 64524 47636 64525 47700
rect 64459 47635 64525 47636
rect 64462 6765 64522 47635
rect 64702 44592 65322 54288
rect 67702 82240 68322 87000
rect 67702 82176 67740 82240
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82176 68322 82240
rect 67702 82160 68322 82176
rect 67702 82096 67740 82160
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82096 68322 82160
rect 67702 82080 68322 82096
rect 67702 82016 67740 82080
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82016 68322 82080
rect 67702 82000 68322 82016
rect 67702 81936 67740 82000
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81936 68322 82000
rect 67702 72240 68322 81936
rect 67702 72176 67740 72240
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72176 68322 72240
rect 67702 72160 68322 72176
rect 67702 72096 67740 72160
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72096 68322 72160
rect 67702 72080 68322 72096
rect 67702 72016 67740 72080
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72016 68322 72080
rect 67702 72000 68322 72016
rect 67702 71936 67740 72000
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71936 68322 72000
rect 67702 62240 68322 71936
rect 67702 62176 67740 62240
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62176 68322 62240
rect 67702 62160 68322 62176
rect 67702 62096 67740 62160
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62096 68322 62160
rect 67702 62080 68322 62096
rect 67702 62016 67740 62080
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62016 68322 62080
rect 67702 62000 68322 62016
rect 67702 61936 67740 62000
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61936 68322 62000
rect 67702 52240 68322 61936
rect 67702 52176 67740 52240
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52176 68322 52240
rect 67702 52160 68322 52176
rect 67702 52096 67740 52160
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52096 68322 52160
rect 67702 52080 68322 52096
rect 67702 52016 67740 52080
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52016 68322 52080
rect 67702 52000 68322 52016
rect 67702 51936 67740 52000
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51936 68322 52000
rect 65563 48108 65629 48109
rect 65563 48044 65564 48108
rect 65628 48044 65629 48108
rect 65563 48043 65629 48044
rect 64702 44528 64740 44592
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 65322 44592
rect 64702 44512 65322 44528
rect 64702 44448 64740 44512
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 65322 44512
rect 64702 44432 65322 44448
rect 64702 44368 64740 44432
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 65322 44432
rect 64702 44352 65322 44368
rect 64702 44288 64740 44352
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 65322 44352
rect 64702 34592 65322 44288
rect 64702 34528 64740 34592
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 65322 34592
rect 64702 34512 65322 34528
rect 64702 34448 64740 34512
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 65322 34512
rect 64702 34432 65322 34448
rect 64702 34368 64740 34432
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 65322 34432
rect 64702 34352 65322 34368
rect 64702 34288 64740 34352
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 65322 34352
rect 64702 24592 65322 34288
rect 64702 24528 64740 24592
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 65322 24592
rect 64702 24512 65322 24528
rect 64702 24448 64740 24512
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 65322 24512
rect 64702 24432 65322 24448
rect 64702 24368 64740 24432
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 65322 24432
rect 64702 24352 65322 24368
rect 64702 24288 64740 24352
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 65322 24352
rect 64702 14592 65322 24288
rect 64702 14528 64740 14592
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 65322 14592
rect 64702 14512 65322 14528
rect 64702 14448 64740 14512
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 65322 14512
rect 64702 14432 65322 14448
rect 64702 14368 64740 14432
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 65322 14432
rect 64702 14352 65322 14368
rect 64702 14288 64740 14352
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 65322 14352
rect 64459 6764 64525 6765
rect 64459 6700 64460 6764
rect 64524 6700 64525 6764
rect 64459 6699 64525 6700
rect 64275 4996 64341 4997
rect 64275 4932 64276 4996
rect 64340 4932 64341 4996
rect 64275 4931 64341 4932
rect 63171 4860 63237 4861
rect 63171 4796 63172 4860
rect 63236 4796 63237 4860
rect 63171 4795 63237 4796
rect 61702 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2176 61900 2240
rect 61964 2176 61980 2240
rect 62044 2176 62060 2240
rect 62124 2176 62140 2240
rect 62204 2176 62220 2240
rect 62284 2176 62322 2240
rect 61702 2160 62322 2176
rect 61702 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2096 61900 2160
rect 61964 2096 61980 2160
rect 62044 2096 62060 2160
rect 62124 2096 62140 2160
rect 62204 2096 62220 2160
rect 62284 2096 62322 2160
rect 61702 2080 62322 2096
rect 61702 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2016 61900 2080
rect 61964 2016 61980 2080
rect 62044 2016 62060 2080
rect 62124 2016 62140 2080
rect 62204 2016 62220 2080
rect 62284 2016 62322 2080
rect 61702 2000 62322 2016
rect 61702 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1936 61900 2000
rect 61964 1936 61980 2000
rect 62044 1936 62060 2000
rect 62124 1936 62140 2000
rect 62204 1936 62220 2000
rect 62284 1936 62322 2000
rect 61702 0 62322 1936
rect 64702 4592 65322 14288
rect 65566 11661 65626 48043
rect 67702 42240 68322 51936
rect 67702 42176 67740 42240
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42176 68322 42240
rect 67702 42160 68322 42176
rect 67702 42096 67740 42160
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42096 68322 42160
rect 67702 42080 68322 42096
rect 67702 42016 67740 42080
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42016 68322 42080
rect 67702 42000 68322 42016
rect 67702 41936 67740 42000
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41936 68322 42000
rect 65747 40900 65813 40901
rect 65747 40836 65748 40900
rect 65812 40836 65813 40900
rect 65747 40835 65813 40836
rect 65563 11660 65629 11661
rect 65563 11596 65564 11660
rect 65628 11596 65629 11660
rect 65563 11595 65629 11596
rect 65563 11524 65629 11525
rect 65563 11460 65564 11524
rect 65628 11460 65629 11524
rect 65563 11459 65629 11460
rect 65566 7717 65626 11459
rect 65563 7716 65629 7717
rect 65563 7652 65564 7716
rect 65628 7652 65629 7716
rect 65563 7651 65629 7652
rect 65750 7581 65810 40835
rect 65931 38724 65997 38725
rect 65931 38660 65932 38724
rect 65996 38660 65997 38724
rect 65931 38659 65997 38660
rect 65747 7580 65813 7581
rect 65747 7516 65748 7580
rect 65812 7516 65813 7580
rect 65747 7515 65813 7516
rect 65934 6221 65994 38659
rect 67702 32240 68322 41936
rect 70702 84592 71322 87000
rect 70702 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84528 71322 84592
rect 70702 84512 71322 84528
rect 70702 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84448 71322 84512
rect 70702 84432 71322 84448
rect 70702 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84368 71322 84432
rect 70702 84352 71322 84368
rect 70702 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84288 71322 84352
rect 70702 74592 71322 84288
rect 70702 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74528 71322 74592
rect 70702 74512 71322 74528
rect 70702 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74448 71322 74512
rect 70702 74432 71322 74448
rect 70702 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74368 71322 74432
rect 70702 74352 71322 74368
rect 70702 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74288 71322 74352
rect 70702 64592 71322 74288
rect 70702 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64528 71322 64592
rect 70702 64512 71322 64528
rect 70702 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64448 71322 64512
rect 70702 64432 71322 64448
rect 70702 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64368 71322 64432
rect 70702 64352 71322 64368
rect 70702 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64288 71322 64352
rect 70702 54592 71322 64288
rect 70702 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54528 71322 54592
rect 70702 54512 71322 54528
rect 70702 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54448 71322 54512
rect 70702 54432 71322 54448
rect 70702 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54368 71322 54432
rect 70702 54352 71322 54368
rect 70702 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54288 71322 54352
rect 70702 44592 71322 54288
rect 70702 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44528 71322 44592
rect 70702 44512 71322 44528
rect 70702 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44448 71322 44512
rect 70702 44432 71322 44448
rect 70702 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44368 71322 44432
rect 70702 44352 71322 44368
rect 70702 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44288 71322 44352
rect 70702 34592 71322 44288
rect 70702 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34528 71322 34592
rect 70702 34512 71322 34528
rect 70702 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34448 71322 34512
rect 70702 34432 71322 34448
rect 70702 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34368 71322 34432
rect 70702 34352 71322 34368
rect 70702 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34288 71322 34352
rect 68507 33284 68573 33285
rect 68507 33220 68508 33284
rect 68572 33220 68573 33284
rect 68507 33219 68573 33220
rect 67702 32176 67740 32240
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32176 68322 32240
rect 67702 32160 68322 32176
rect 67702 32096 67740 32160
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32096 68322 32160
rect 67702 32080 68322 32096
rect 67702 32016 67740 32080
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32016 68322 32080
rect 67702 32000 68322 32016
rect 67702 31936 67740 32000
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31936 68322 32000
rect 66299 23492 66365 23493
rect 66299 23428 66300 23492
rect 66364 23428 66365 23492
rect 66299 23427 66365 23428
rect 66483 23492 66549 23493
rect 66483 23428 66484 23492
rect 66548 23428 66549 23492
rect 66483 23427 66549 23428
rect 66115 11660 66181 11661
rect 66115 11596 66116 11660
rect 66180 11596 66181 11660
rect 66115 11595 66181 11596
rect 65931 6220 65997 6221
rect 65931 6156 65932 6220
rect 65996 6156 65997 6220
rect 65931 6155 65997 6156
rect 64702 4528 64740 4592
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 65322 4592
rect 64702 4512 65322 4528
rect 64702 4448 64740 4512
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 65322 4512
rect 64702 4432 65322 4448
rect 64702 4368 64740 4432
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 65322 4432
rect 64702 4352 65322 4368
rect 64702 4288 64740 4352
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 65322 4352
rect 64702 0 65322 4288
rect 66118 4045 66178 11595
rect 66115 4044 66181 4045
rect 66115 3980 66116 4044
rect 66180 3980 66181 4044
rect 66115 3979 66181 3980
rect 66302 3365 66362 23427
rect 66486 5269 66546 23427
rect 67702 22240 68322 31936
rect 67702 22176 67740 22240
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22176 68322 22240
rect 67702 22160 68322 22176
rect 67702 22096 67740 22160
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22096 68322 22160
rect 67702 22080 68322 22096
rect 67702 22016 67740 22080
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22016 68322 22080
rect 67702 22000 68322 22016
rect 67702 21936 67740 22000
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21936 68322 22000
rect 66667 19140 66733 19141
rect 66667 19076 66668 19140
rect 66732 19076 66733 19140
rect 66667 19075 66733 19076
rect 66670 6901 66730 19075
rect 67702 12240 68322 21936
rect 67702 12176 67740 12240
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12176 68322 12240
rect 67702 12160 68322 12176
rect 67702 12096 67740 12160
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12096 68322 12160
rect 67702 12080 68322 12096
rect 67702 12016 67740 12080
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12016 68322 12080
rect 67702 12000 68322 12016
rect 67702 11936 67740 12000
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11936 68322 12000
rect 66667 6900 66733 6901
rect 66667 6836 66668 6900
rect 66732 6836 66733 6900
rect 66667 6835 66733 6836
rect 66483 5268 66549 5269
rect 66483 5204 66484 5268
rect 66548 5204 66549 5268
rect 66483 5203 66549 5204
rect 66299 3364 66365 3365
rect 66299 3300 66300 3364
rect 66364 3300 66365 3364
rect 66299 3299 66365 3300
rect 67702 2240 68322 11936
rect 68510 5677 68570 33219
rect 70702 24592 71322 34288
rect 70702 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24528 71322 24592
rect 70702 24512 71322 24528
rect 70702 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24448 71322 24512
rect 70702 24432 71322 24448
rect 70702 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24368 71322 24432
rect 70702 24352 71322 24368
rect 70702 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24288 71322 24352
rect 70702 14592 71322 24288
rect 70702 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14528 71322 14592
rect 70702 14512 71322 14528
rect 70702 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14448 71322 14512
rect 70702 14432 71322 14448
rect 70702 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14368 71322 14432
rect 70702 14352 71322 14368
rect 70702 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14288 71322 14352
rect 68507 5676 68573 5677
rect 68507 5612 68508 5676
rect 68572 5612 68573 5676
rect 68507 5611 68573 5612
rect 67702 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2176 68322 2240
rect 67702 2160 68322 2176
rect 67702 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2096 68322 2160
rect 67702 2080 68322 2096
rect 67702 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2016 68322 2080
rect 67702 2000 68322 2016
rect 67702 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1936 68322 2000
rect 67702 0 68322 1936
rect 70702 4592 71322 14288
rect 70702 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4528 71322 4592
rect 70702 4512 71322 4528
rect 70702 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4448 71322 4512
rect 70702 4432 71322 4448
rect 70702 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4368 71322 4432
rect 70702 4352 71322 4368
rect 70702 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4288 71322 4352
rect 70702 0 71322 4288
rect 73702 82240 74322 87000
rect 73702 82176 73740 82240
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 74322 82240
rect 73702 82160 74322 82176
rect 73702 82096 73740 82160
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 74322 82160
rect 73702 82080 74322 82096
rect 73702 82016 73740 82080
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 74322 82080
rect 73702 82000 74322 82016
rect 73702 81936 73740 82000
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 74322 82000
rect 73702 72240 74322 81936
rect 73702 72176 73740 72240
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 74322 72240
rect 73702 72160 74322 72176
rect 73702 72096 73740 72160
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 74322 72160
rect 73702 72080 74322 72096
rect 73702 72016 73740 72080
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 74322 72080
rect 73702 72000 74322 72016
rect 73702 71936 73740 72000
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 74322 72000
rect 73702 62240 74322 71936
rect 73702 62176 73740 62240
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 74322 62240
rect 73702 62160 74322 62176
rect 73702 62096 73740 62160
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 74322 62160
rect 73702 62080 74322 62096
rect 73702 62016 73740 62080
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 74322 62080
rect 73702 62000 74322 62016
rect 73702 61936 73740 62000
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 74322 62000
rect 73702 52240 74322 61936
rect 73702 52176 73740 52240
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 74322 52240
rect 73702 52160 74322 52176
rect 73702 52096 73740 52160
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 74322 52160
rect 73702 52080 74322 52096
rect 73702 52016 73740 52080
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 74322 52080
rect 73702 52000 74322 52016
rect 73702 51936 73740 52000
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 74322 52000
rect 73702 42240 74322 51936
rect 73702 42176 73740 42240
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 74322 42240
rect 73702 42160 74322 42176
rect 73702 42096 73740 42160
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 74322 42160
rect 73702 42080 74322 42096
rect 73702 42016 73740 42080
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 74322 42080
rect 73702 42000 74322 42016
rect 73702 41936 73740 42000
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 74322 42000
rect 73702 32240 74322 41936
rect 73702 32176 73740 32240
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 74322 32240
rect 73702 32160 74322 32176
rect 73702 32096 73740 32160
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 74322 32160
rect 73702 32080 74322 32096
rect 73702 32016 73740 32080
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 74322 32080
rect 73702 32000 74322 32016
rect 73702 31936 73740 32000
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 74322 32000
rect 73702 22240 74322 31936
rect 73702 22176 73740 22240
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 74322 22240
rect 73702 22160 74322 22176
rect 73702 22096 73740 22160
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 74322 22160
rect 73702 22080 74322 22096
rect 73702 22016 73740 22080
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 74322 22080
rect 73702 22000 74322 22016
rect 73702 21936 73740 22000
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 74322 22000
rect 73702 12240 74322 21936
rect 73702 12176 73740 12240
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 74322 12240
rect 73702 12160 74322 12176
rect 73702 12096 73740 12160
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 74322 12160
rect 73702 12080 74322 12096
rect 73702 12016 73740 12080
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 74322 12080
rect 73702 12000 74322 12016
rect 73702 11936 73740 12000
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 74322 12000
rect 73702 2240 74322 11936
rect 73702 2176 73740 2240
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 74322 2240
rect 73702 2160 74322 2176
rect 73702 2096 73740 2160
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 74322 2160
rect 73702 2080 74322 2096
rect 73702 2016 73740 2080
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 74322 2080
rect 73702 2000 74322 2016
rect 73702 1936 73740 2000
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 74322 2000
rect 73702 0 74322 1936
use sky130_fd_sc_hd__nor2b_4  _049_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 44436 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _050_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _051_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 30912 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25944 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _053_
timestamp 1704896540
transform -1 0 30360 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1704896540
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _055_
timestamp 1704896540
transform -1 0 29808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp 1704896540
transform -1 0 26772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _057_
timestamp 1704896540
transform -1 0 29164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp 1704896540
transform -1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _059_
timestamp 1704896540
transform -1 0 28520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp 1704896540
transform -1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _061_
timestamp 1704896540
transform 1 0 27048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp 1704896540
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _063_
timestamp 1704896540
transform 1 0 26312 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp 1704896540
transform 1 0 29440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _065_
timestamp 1704896540
transform 1 0 25852 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp 1704896540
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _067_
timestamp 1704896540
transform 1 0 24196 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp 1704896540
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _069_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 35052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _070_
timestamp 1704896540
transform 1 0 25392 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp 1704896540
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _072_
timestamp 1704896540
transform 1 0 24748 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _073_
timestamp 1704896540
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _074_
timestamp 1704896540
transform 1 0 24288 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp 1704896540
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _076_
timestamp 1704896540
transform 1 0 23276 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp 1704896540
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _078_
timestamp 1704896540
transform 1 0 23736 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp 1704896540
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _080_
timestamp 1704896540
transform 1 0 25760 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp 1704896540
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _082_
timestamp 1704896540
transform 1 0 27508 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp 1704896540
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _084_
timestamp 1704896540
transform 1 0 44068 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp 1704896540
transform 1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _086_
timestamp 1704896540
transform 1 0 46092 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp 1704896540
transform 1 0 47472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _088_
timestamp 1704896540
transform 1 0 46644 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp 1704896540
transform 1 0 49036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1704896540
transform -1 0 61364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1704896540
transform -1 0 53360 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp 1704896540
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _093_
timestamp 1704896540
transform -1 0 55016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp 1704896540
transform 1 0 54648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _095_
timestamp 1704896540
transform -1 0 56580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp 1704896540
transform 1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _097_
timestamp 1704896540
transform -1 0 58236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp 1704896540
transform 1 0 57776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _099_
timestamp 1704896540
transform -1 0 59800 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp 1704896540
transform 1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _101_
timestamp 1704896540
transform -1 0 61732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp 1704896540
transform 1 0 61180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _103_
timestamp 1704896540
transform 1 0 62928 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp 1704896540
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _105_
timestamp 1704896540
transform -1 0 65136 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _106_
timestamp 1704896540
transform -1 0 64860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _107_
timestamp 1704896540
transform 1 0 66148 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1704896540
transform -1 0 66516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _109_
timestamp 1704896540
transform -1 0 68540 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _110_
timestamp 1704896540
transform 1 0 68080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _111_
timestamp 1704896540
transform -1 0 70472 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1704896540
transform -1 0 69920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _113_
timestamp 1704896540
transform -1 0 71944 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1704896540
transform -1 0 71484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _115_
timestamp 1704896540
transform -1 0 73692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _116_
timestamp 1704896540
transform 1 0 72864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _117_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 30728 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _118_
timestamp 1704896540
transform -1 0 23736 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1704896540
transform -1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25852 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _122_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20608 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20056 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 40388 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1704896540
transform -1 0 37076 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1704896540
transform 1 0 65596 0 1 33728
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2392 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6256 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7360 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8464 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8832 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9936 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11408 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12512 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13984 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_159
timestamp 1704896540
transform 1 0 15640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1704896540
transform 1 0 18952 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_220 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21252 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21712 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1704896540
transform 1 0 24288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_337
timestamp 1704896540
transform 1 0 32016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1704896540
transform 1 0 34592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_393
timestamp 1704896540
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39468 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1704896540
transform 1 0 41952 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1704896540
transform 1 0 49680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1704896540
transform 1 0 52256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1704896540
transform 1 0 54832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1704896540
transform 1 0 57408 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_617
timestamp 1704896540
transform 1 0 57776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_642
timestamp 1704896540
transform 1 0 60076 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1704896540
transform 1 0 62560 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1704896540
transform 1 0 65136 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_707
timestamp 1704896540
transform 1 0 66056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_724
timestamp 1704896540
transform 1 0 67620 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_753
timestamp 1704896540
transform 1 0 70288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_757
timestamp 1704896540
transform 1 0 70656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_761
timestamp 1704896540
transform 1 0 71024 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1288 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2392 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3496 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4600 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6256 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7360 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8464 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9568 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10672 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11224 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11408 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12512 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13616 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14720 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15824 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16560 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21528 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_271
timestamp 1704896540
transform 1 0 25944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_297
timestamp 1704896540
transform 1 0 28336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_337
timestamp 1704896540
transform 1 0 32016 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1704896540
transform 1 0 32384 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1704896540
transform 1 0 36892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_393
timestamp 1704896540
transform 1 0 37168 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_410
timestamp 1704896540
transform 1 0 38732 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_430
timestamp 1704896540
transform 1 0 40572 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_434
timestamp 1704896540
transform 1 0 40940 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1704896540
transform 1 0 42136 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_449
timestamp 1704896540
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_454
timestamp 1704896540
transform 1 0 42780 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1704896540
transform 1 0 47288 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_505
timestamp 1704896540
transform 1 0 47472 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_509
timestamp 1704896540
transform 1 0 47840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_540
timestamp 1704896540
transform 1 0 50692 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_544
timestamp 1704896540
transform 1 0 51060 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1704896540
transform 1 0 52440 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_561
timestamp 1704896540
transform 1 0 52624 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_588
timestamp 1704896540
transform 1 0 55108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_631
timestamp 1704896540
transform 1 0 59064 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_670
timestamp 1704896540
transform 1 0 62652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_681
timestamp 1704896540
transform 1 0 63664 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_737
timestamp 1704896540
transform 1 0 68816 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_774
timestamp 1704896540
transform 1 0 72220 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_783
timestamp 1704896540
transform 1 0 73048 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_793
timestamp 1704896540
transform 1 0 73968 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3496 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8648 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 11040 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13800 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15088 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_173
timestamp 1704896540
transform 1 0 16928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 1704896540
transform 1 0 24288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_296
timestamp 1704896540
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_317
timestamp 1704896540
transform 1 0 30176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_350
timestamp 1704896540
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1704896540
transform 1 0 34316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_365
timestamp 1704896540
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_388
timestamp 1704896540
transform 1 0 36708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_400
timestamp 1704896540
transform 1 0 37812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_412
timestamp 1704896540
transform 1 0 38916 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1704896540
transform 1 0 39744 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1704896540
transform 1 0 40848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_445
timestamp 1704896540
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_449
timestamp 1704896540
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_458
timestamp 1704896540
transform 1 0 43148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_485
timestamp 1704896540
transform 1 0 45632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_489
timestamp 1704896540
transform 1 0 46000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_512
timestamp 1704896540
transform 1 0 48116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_520
timestamp 1704896540
transform 1 0 48852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_530
timestamp 1704896540
transform 1 0 49772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1704896540
transform 1 0 50048 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1704896540
transform 1 0 51152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_557
timestamp 1704896540
transform 1 0 52256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_565
timestamp 1704896540
transform 1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_576
timestamp 1704896540
transform 1 0 54004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_585
timestamp 1704896540
transform 1 0 54832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_601
timestamp 1704896540
transform 1 0 56304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_609
timestamp 1704896540
transform 1 0 57040 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_620
timestamp 1704896540
transform 1 0 58052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_632
timestamp 1704896540
transform 1 0 59156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_645
timestamp 1704896540
transform 1 0 60352 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_654
timestamp 1704896540
transform 1 0 61180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_680
timestamp 1704896540
transform 1 0 63572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_692
timestamp 1704896540
transform 1 0 64676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_701
timestamp 1704896540
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_710
timestamp 1704896540
transform 1 0 66332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_718
timestamp 1704896540
transform 1 0 67068 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_726
timestamp 1704896540
transform 1 0 67804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_738
timestamp 1704896540
transform 1 0 68908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_750
timestamp 1704896540
transform 1 0 70012 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_765
timestamp 1704896540
transform 1 0 71392 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_777
timestamp 1704896540
transform 1 0 72496 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_789
timestamp 1704896540
transform 1 0 73600 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16376 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_187
timestamp 1704896540
transform 1 0 18216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_249
timestamp 1704896540
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_261
timestamp 1704896540
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_274
timestamp 1704896540
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_295
timestamp 1704896540
transform 1 0 28152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_326
timestamp 1704896540
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 1704896540
transform 1 0 31740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_349
timestamp 1704896540
transform 1 0 33120 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_366
timestamp 1704896540
transform 1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_385
timestamp 1704896540
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1704896540
transform 1 0 37168 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1704896540
transform 1 0 38272 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1704896540
transform 1 0 39376 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1704896540
transform 1 0 40480 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1704896540
transform 1 0 41584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1704896540
transform 1 0 42136 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1704896540
transform 1 0 42320 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1704896540
transform 1 0 43424 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1704896540
transform 1 0 44528 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_485
timestamp 1704896540
transform 1 0 45632 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_491
timestamp 1704896540
transform 1 0 46184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1704896540
transform 1 0 47288 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_508
timestamp 1704896540
transform 1 0 47748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_520
timestamp 1704896540
transform 1 0 48852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_525
timestamp 1704896540
transform 1 0 49312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_537
timestamp 1704896540
transform 1 0 50416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_549
timestamp 1704896540
transform 1 0 51520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_557
timestamp 1704896540
transform 1 0 52256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_561
timestamp 1704896540
transform 1 0 52624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_567
timestamp 1704896540
transform 1 0 53176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_575
timestamp 1704896540
transform 1 0 53912 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_586
timestamp 1704896540
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_598
timestamp 1704896540
transform 1 0 56028 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_603
timestamp 1704896540
transform 1 0 56488 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1704896540
transform 1 0 57592 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_620
timestamp 1704896540
transform 1 0 58052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_632
timestamp 1704896540
transform 1 0 59156 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_638
timestamp 1704896540
transform 1 0 59708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_650
timestamp 1704896540
transform 1 0 60812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_657
timestamp 1704896540
transform 1 0 61456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_669
timestamp 1704896540
transform 1 0 62560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_673
timestamp 1704896540
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_677
timestamp 1704896540
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_689
timestamp 1704896540
transform 1 0 64400 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_694
timestamp 1704896540
transform 1 0 64860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_706
timestamp 1704896540
transform 1 0 65964 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_712
timestamp 1704896540
transform 1 0 66516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_724
timestamp 1704896540
transform 1 0 67620 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_732
timestamp 1704896540
transform 1 0 68356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_744
timestamp 1704896540
transform 1 0 69460 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_749
timestamp 1704896540
transform 1 0 69920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_761
timestamp 1704896540
transform 1 0 71024 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_766
timestamp 1704896540
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_778
timestamp 1704896540
transform 1 0 72588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1704896540
transform 1 0 73232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_797
timestamp 1704896540
transform 1 0 74336 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8648 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9936 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15088 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18952 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_217
timestamp 1704896540
transform 1 0 20976 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_229
timestamp 1704896540
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_233
timestamp 1704896540
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 1704896540
transform 1 0 23736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1704896540
transform 1 0 24104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_253
timestamp 1704896540
transform 1 0 24288 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_257
timestamp 1704896540
transform 1 0 24656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_275
timestamp 1704896540
transform 1 0 26312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_283
timestamp 1704896540
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_295
timestamp 1704896540
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1704896540
transform 1 0 29256 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1704896540
transform 1 0 29440 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_321
timestamp 1704896540
transform 1 0 30544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_327
timestamp 1704896540
transform 1 0 31096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_331
timestamp 1704896540
transform 1 0 31464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_336
timestamp 1704896540
transform 1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_342
timestamp 1704896540
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_349
timestamp 1704896540
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_361
timestamp 1704896540
transform 1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1704896540
transform 1 0 34592 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1704896540
transform 1 0 35696 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1704896540
transform 1 0 36800 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1704896540
transform 1 0 37904 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1704896540
transform 1 0 39008 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1704896540
transform 1 0 39560 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1704896540
transform 1 0 39744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1704896540
transform 1 0 40848 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1704896540
transform 1 0 41952 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1704896540
transform 1 0 43056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1704896540
transform 1 0 44160 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1704896540
transform 1 0 44712 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1704896540
transform 1 0 44896 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1704896540
transform 1 0 46000 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1704896540
transform 1 0 47104 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1704896540
transform 1 0 48208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 1704896540
transform 1 0 49312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1704896540
transform 1 0 49864 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1704896540
transform 1 0 50048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1704896540
transform 1 0 51152 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1704896540
transform 1 0 52256 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1704896540
transform 1 0 53360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1704896540
transform 1 0 54464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1704896540
transform 1 0 55016 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1704896540
transform 1 0 55200 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1704896540
transform 1 0 56304 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1704896540
transform 1 0 57408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1704896540
transform 1 0 58512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1704896540
transform 1 0 59616 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1704896540
transform 1 0 60168 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1704896540
transform 1 0 60352 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1704896540
transform 1 0 61456 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1704896540
transform 1 0 62560 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1704896540
transform 1 0 63664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1704896540
transform 1 0 64768 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1704896540
transform 1 0 65320 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1704896540
transform 1 0 65504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1704896540
transform 1 0 66608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_725
timestamp 1704896540
transform 1 0 67712 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_737
timestamp 1704896540
transform 1 0 68816 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_749
timestamp 1704896540
transform 1 0 69920 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_755
timestamp 1704896540
transform 1 0 70472 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1704896540
transform 1 0 70656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1704896540
transform 1 0 71760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1704896540
transform 1 0 72864 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_793
timestamp 1704896540
transform 1 0 73968 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6072 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10672 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11224 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13616 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16376 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_197
timestamp 1704896540
transform 1 0 19136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_204
timestamp 1704896540
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_216
timestamp 1704896540
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22816 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1704896540
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1704896540
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 26128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_287
timestamp 1704896540
transform 1 0 27416 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_294
timestamp 1704896540
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_306
timestamp 1704896540
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_320
timestamp 1704896540
transform 1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_330
timestamp 1704896540
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1704896540
transform 1 0 32016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1704896540
transform 1 0 33120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_361
timestamp 1704896540
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_365
timestamp 1704896540
transform 1 0 34592 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_370
timestamp 1704896540
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_382
timestamp 1704896540
transform 1 0 36156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1704896540
transform 1 0 36892 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1704896540
transform 1 0 37168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1704896540
transform 1 0 38272 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1704896540
transform 1 0 39376 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1704896540
transform 1 0 40480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1704896540
transform 1 0 41584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1704896540
transform 1 0 42136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1704896540
transform 1 0 42320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1704896540
transform 1 0 43424 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1704896540
transform 1 0 44528 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1704896540
transform 1 0 45632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 1704896540
transform 1 0 46736 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1704896540
transform 1 0 47288 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1704896540
transform 1 0 47472 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1704896540
transform 1 0 48576 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1704896540
transform 1 0 49680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1704896540
transform 1 0 50784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 1704896540
transform 1 0 51888 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1704896540
transform 1 0 52440 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1704896540
transform 1 0 52624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1704896540
transform 1 0 53728 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1704896540
transform 1 0 54832 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1704896540
transform 1 0 55936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1704896540
transform 1 0 57040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1704896540
transform 1 0 57592 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1704896540
transform 1 0 57776 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1704896540
transform 1 0 58880 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1704896540
transform 1 0 59984 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1704896540
transform 1 0 61088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1704896540
transform 1 0 62192 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1704896540
transform 1 0 62744 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1704896540
transform 1 0 62928 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1704896540
transform 1 0 64032 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1704896540
transform 1 0 65136 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1704896540
transform 1 0 66240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1704896540
transform 1 0 67344 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1704896540
transform 1 0 67896 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1704896540
transform 1 0 68080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1704896540
transform 1 0 69184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1704896540
transform 1 0 70288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1704896540
transform 1 0 71392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1704896540
transform 1 0 72496 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1704896540
transform 1 0 73048 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1704896540
transform 1 0 73232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_797
timestamp 1704896540
transform 1 0 74336 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8096 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8648 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9936 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13800 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15088 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23552 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 24104 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1704896540
transform 1 0 24288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1704896540
transform 1 0 25392 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1704896540
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1704896540
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1704896540
transform 1 0 28704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1704896540
transform 1 0 29256 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1704896540
transform 1 0 29440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1704896540
transform 1 0 30544 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1704896540
transform 1 0 31648 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1704896540
transform 1 0 32752 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_357
timestamp 1704896540
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1704896540
transform 1 0 34592 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1704896540
transform 1 0 35696 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1704896540
transform 1 0 36800 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1704896540
transform 1 0 37904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1704896540
transform 1 0 39008 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1704896540
transform 1 0 39560 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1704896540
transform 1 0 39744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_433
timestamp 1704896540
transform 1 0 40848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_453
timestamp 1704896540
transform 1 0 42688 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_459
timestamp 1704896540
transform 1 0 43240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_473
timestamp 1704896540
transform 1 0 44528 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1704896540
transform 1 0 44896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_489
timestamp 1704896540
transform 1 0 46000 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_495
timestamp 1704896540
transform 1 0 46552 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1704896540
transform 1 0 47104 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1704896540
transform 1 0 48208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 1704896540
transform 1 0 49312 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 1704896540
transform 1 0 49864 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1704896540
transform 1 0 50048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1704896540
transform 1 0 51152 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1704896540
transform 1 0 52256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1704896540
transform 1 0 53360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1704896540
transform 1 0 54464 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1704896540
transform 1 0 55016 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1704896540
transform 1 0 55200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1704896540
transform 1 0 56304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1704896540
transform 1 0 57408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1704896540
transform 1 0 58512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1704896540
transform 1 0 59616 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1704896540
transform 1 0 60168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_645
timestamp 1704896540
transform 1 0 60352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_651
timestamp 1704896540
transform 1 0 60904 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_656
timestamp 1704896540
transform 1 0 61364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_668
timestamp 1704896540
transform 1 0 62468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_680
timestamp 1704896540
transform 1 0 63572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_692
timestamp 1704896540
transform 1 0 64676 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1704896540
transform 1 0 65504 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1704896540
transform 1 0 66608 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1704896540
transform 1 0 67712 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1704896540
transform 1 0 68816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1704896540
transform 1 0 69920 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1704896540
transform 1 0 70472 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1704896540
transform 1 0 70656 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1704896540
transform 1 0 71760 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1704896540
transform 1 0 72864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_793
timestamp 1704896540
transform 1 0 73968 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10672 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11224 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16376 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1704896540
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1704896540
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22816 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp 1704896540
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_260
timestamp 1704896540
transform 1 0 24932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_264
timestamp 1704896540
transform 1 0 25300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_293
timestamp 1704896540
transform 1 0 27968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_299
timestamp 1704896540
transform 1 0 28520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_306
timestamp 1704896540
transform 1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_313
timestamp 1704896540
transform 1 0 29808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_319
timestamp 1704896540
transform 1 0 30360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_325
timestamp 1704896540
transform 1 0 30912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_333
timestamp 1704896540
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1704896540
transform 1 0 32016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1704896540
transform 1 0 33120 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1704896540
transform 1 0 34224 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1704896540
transform 1 0 35328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1704896540
transform 1 0 36432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1704896540
transform 1 0 36984 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1704896540
transform 1 0 37168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1704896540
transform 1 0 38272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_417
timestamp 1704896540
transform 1 0 39376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_425
timestamp 1704896540
transform 1 0 40112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_436
timestamp 1704896540
transform 1 0 41124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_449
timestamp 1704896540
transform 1 0 42320 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_455
timestamp 1704896540
transform 1 0 42872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_480
timestamp 1704896540
transform 1 0 45172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 1704896540
transform 1 0 47288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_513
timestamp 1704896540
transform 1 0 48208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_521
timestamp 1704896540
transform 1 0 48944 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_531
timestamp 1704896540
transform 1 0 49864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_543
timestamp 1704896540
transform 1 0 50968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_555
timestamp 1704896540
transform 1 0 52072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 1704896540
transform 1 0 52440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_561
timestamp 1704896540
transform 1 0 52624 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_569
timestamp 1704896540
transform 1 0 53360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_581
timestamp 1704896540
transform 1 0 54464 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_587
timestamp 1704896540
transform 1 0 55016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_599
timestamp 1704896540
transform 1 0 56120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_611
timestamp 1704896540
transform 1 0 57224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1704896540
transform 1 0 57592 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1704896540
transform 1 0 57776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1704896540
transform 1 0 58880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1704896540
transform 1 0 59984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1704896540
transform 1 0 61088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1704896540
transform 1 0 62192 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1704896540
transform 1 0 62744 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1704896540
transform 1 0 62928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1704896540
transform 1 0 64032 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1704896540
transform 1 0 65136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1704896540
transform 1 0 66240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1704896540
transform 1 0 67344 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1704896540
transform 1 0 67896 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1704896540
transform 1 0 68080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_741
timestamp 1704896540
transform 1 0 69184 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_749
timestamp 1704896540
transform 1 0 69920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_755
timestamp 1704896540
transform 1 0 70472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_763
timestamp 1704896540
transform 1 0 71208 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_771
timestamp 1704896540
transform 1 0 71944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1704896540
transform 1 0 73048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_790
timestamp 1704896540
transform 1 0 73692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_798
timestamp 1704896540
transform 1 0 74428 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1704896540
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1704896540
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1704896540
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_113
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1704896540
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1704896540
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_169
timestamp 1704896540
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_181
timestamp 1704896540
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1704896540
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 20240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_221
timestamp 1704896540
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_225
timestamp 1704896540
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_237
timestamp 1704896540
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_241
timestamp 1704896540
transform 1 0 23184 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_263
timestamp 1704896540
transform 1 0 25208 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_274
timestamp 1704896540
transform 1 0 26220 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_281
timestamp 1704896540
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_293
timestamp 1704896540
transform 1 0 27968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 1704896540
transform 1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1704896540
transform 1 0 29440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1704896540
transform 1 0 30544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_333
timestamp 1704896540
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_337
timestamp 1704896540
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_349
timestamp 1704896540
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1704896540
transform 1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_365
timestamp 1704896540
transform 1 0 34592 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_371
timestamp 1704896540
transform 1 0 35144 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_393
timestamp 1704896540
transform 1 0 37168 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_405
timestamp 1704896540
transform 1 0 38272 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_417
timestamp 1704896540
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_421
timestamp 1704896540
transform 1 0 39744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_427
timestamp 1704896540
transform 1 0 40296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1704896540
transform 1 0 44528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_501
timestamp 1704896540
transform 1 0 47104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_529
timestamp 1704896540
transform 1 0 49680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_533
timestamp 1704896540
transform 1 0 50048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_545
timestamp 1704896540
transform 1 0 51152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_554
timestamp 1704896540
transform 1 0 51980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_585
timestamp 1704896540
transform 1 0 54832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_597
timestamp 1704896540
transform 1 0 55936 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_604
timestamp 1704896540
transform 1 0 56580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_622
timestamp 1704896540
transform 1 0 58236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_639
timestamp 1704896540
transform 1 0 59800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1704896540
transform 1 0 60168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_645
timestamp 1704896540
transform 1 0 60352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_653
timestamp 1704896540
transform 1 0 61088 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_660
timestamp 1704896540
transform 1 0 61732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_678
timestamp 1704896540
transform 1 0 63388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_690
timestamp 1704896540
transform 1 0 64492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_697
timestamp 1704896540
transform 1 0 65136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_701
timestamp 1704896540
transform 1 0 65504 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_707
timestamp 1704896540
transform 1 0 66056 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1704896540
transform 1 0 66608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_725
timestamp 1704896540
transform 1 0 67712 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_734
timestamp 1704896540
transform 1 0 68540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_746
timestamp 1704896540
transform 1 0 69644 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_754
timestamp 1704896540
transform 1 0 70380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1704896540
transform 1 0 70656 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1704896540
transform 1 0 71760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_781
timestamp 1704896540
transform 1 0 72864 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_785
timestamp 1704896540
transform 1 0 73232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_797
timestamp 1704896540
transform 1 0 74336 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_702
timestamp 1704896540
transform 1 0 65596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_714
timestamp 1704896540
transform 1 0 66700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_726
timestamp 1704896540
transform 1 0 67804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_738
timestamp 1704896540
transform 1 0 68908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_750
timestamp 1704896540
transform 1 0 70012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_754
timestamp 1704896540
transform 1 0 70380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_756
timestamp 1704896540
transform 1 0 70564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_768
timestamp 1704896540
transform 1 0 71668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_780
timestamp 1704896540
transform 1 0 72772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_792
timestamp 1704896540
transform 1 0 73876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_800
timestamp 1704896540
transform 1 0 74612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_702
timestamp 1704896540
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_714
timestamp 1704896540
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_726
timestamp 1704896540
transform 1 0 67804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_728
timestamp 1704896540
transform 1 0 67988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_740
timestamp 1704896540
transform 1 0 69092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_752
timestamp 1704896540
transform 1 0 70196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_764
timestamp 1704896540
transform 1 0 71300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_776
timestamp 1704896540
transform 1 0 72404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_782
timestamp 1704896540
transform 1 0 72956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_784
timestamp 1704896540
transform 1 0 73140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_796
timestamp 1704896540
transform 1 0 74244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_800
timestamp 1704896540
transform 1 0 74612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_702
timestamp 1704896540
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_714
timestamp 1704896540
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_726
timestamp 1704896540
transform 1 0 67804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_738
timestamp 1704896540
transform 1 0 68908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_750
timestamp 1704896540
transform 1 0 70012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_754
timestamp 1704896540
transform 1 0 70380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_756
timestamp 1704896540
transform 1 0 70564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_768
timestamp 1704896540
transform 1 0 71668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_780
timestamp 1704896540
transform 1 0 72772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_792
timestamp 1704896540
transform 1 0 73876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_800
timestamp 1704896540
transform 1 0 74612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_702
timestamp 1704896540
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_714
timestamp 1704896540
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_726
timestamp 1704896540
transform 1 0 67804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_728
timestamp 1704896540
transform 1 0 67988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_740
timestamp 1704896540
transform 1 0 69092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_752
timestamp 1704896540
transform 1 0 70196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_764
timestamp 1704896540
transform 1 0 71300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_776
timestamp 1704896540
transform 1 0 72404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_782
timestamp 1704896540
transform 1 0 72956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_784
timestamp 1704896540
transform 1 0 73140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_796
timestamp 1704896540
transform 1 0 74244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_800
timestamp 1704896540
transform 1 0 74612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_702
timestamp 1704896540
transform 1 0 65596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_714
timestamp 1704896540
transform 1 0 66700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_726
timestamp 1704896540
transform 1 0 67804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_738
timestamp 1704896540
transform 1 0 68908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_750
timestamp 1704896540
transform 1 0 70012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_754
timestamp 1704896540
transform 1 0 70380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_756
timestamp 1704896540
transform 1 0 70564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_768
timestamp 1704896540
transform 1 0 71668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_780
timestamp 1704896540
transform 1 0 72772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_792
timestamp 1704896540
transform 1 0 73876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_800
timestamp 1704896540
transform 1 0 74612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_702
timestamp 1704896540
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_714
timestamp 1704896540
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_726
timestamp 1704896540
transform 1 0 67804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_728
timestamp 1704896540
transform 1 0 67988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_740
timestamp 1704896540
transform 1 0 69092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_752
timestamp 1704896540
transform 1 0 70196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_764
timestamp 1704896540
transform 1 0 71300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_776
timestamp 1704896540
transform 1 0 72404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_782
timestamp 1704896540
transform 1 0 72956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_784
timestamp 1704896540
transform 1 0 73140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_796
timestamp 1704896540
transform 1 0 74244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_800
timestamp 1704896540
transform 1 0 74612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_702
timestamp 1704896540
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_714
timestamp 1704896540
transform 1 0 66700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_726
timestamp 1704896540
transform 1 0 67804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_738
timestamp 1704896540
transform 1 0 68908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_750
timestamp 1704896540
transform 1 0 70012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_754
timestamp 1704896540
transform 1 0 70380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_756
timestamp 1704896540
transform 1 0 70564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_768
timestamp 1704896540
transform 1 0 71668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_780
timestamp 1704896540
transform 1 0 72772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_792
timestamp 1704896540
transform 1 0 73876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_800
timestamp 1704896540
transform 1 0 74612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_702
timestamp 1704896540
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_714
timestamp 1704896540
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_726
timestamp 1704896540
transform 1 0 67804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_728
timestamp 1704896540
transform 1 0 67988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_740
timestamp 1704896540
transform 1 0 69092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_752
timestamp 1704896540
transform 1 0 70196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_764
timestamp 1704896540
transform 1 0 71300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_776
timestamp 1704896540
transform 1 0 72404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_782
timestamp 1704896540
transform 1 0 72956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_784
timestamp 1704896540
transform 1 0 73140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_796
timestamp 1704896540
transform 1 0 74244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_800
timestamp 1704896540
transform 1 0 74612 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_702
timestamp 1704896540
transform 1 0 65596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_714
timestamp 1704896540
transform 1 0 66700 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_726
timestamp 1704896540
transform 1 0 67804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_738
timestamp 1704896540
transform 1 0 68908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_750
timestamp 1704896540
transform 1 0 70012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_754
timestamp 1704896540
transform 1 0 70380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_756
timestamp 1704896540
transform 1 0 70564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_768
timestamp 1704896540
transform 1 0 71668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_780
timestamp 1704896540
transform 1 0 72772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_792
timestamp 1704896540
transform 1 0 73876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_800
timestamp 1704896540
transform 1 0 74612 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_702
timestamp 1704896540
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_714
timestamp 1704896540
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_726
timestamp 1704896540
transform 1 0 67804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_728
timestamp 1704896540
transform 1 0 67988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_740
timestamp 1704896540
transform 1 0 69092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_752
timestamp 1704896540
transform 1 0 70196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_764
timestamp 1704896540
transform 1 0 71300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_776
timestamp 1704896540
transform 1 0 72404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_782
timestamp 1704896540
transform 1 0 72956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_784
timestamp 1704896540
transform 1 0 73140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_796
timestamp 1704896540
transform 1 0 74244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_800
timestamp 1704896540
transform 1 0 74612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_702
timestamp 1704896540
transform 1 0 65596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_714
timestamp 1704896540
transform 1 0 66700 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_726
timestamp 1704896540
transform 1 0 67804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_738
timestamp 1704896540
transform 1 0 68908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_750
timestamp 1704896540
transform 1 0 70012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_754
timestamp 1704896540
transform 1 0 70380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_756
timestamp 1704896540
transform 1 0 70564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_768
timestamp 1704896540
transform 1 0 71668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_780
timestamp 1704896540
transform 1 0 72772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_792
timestamp 1704896540
transform 1 0 73876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_800
timestamp 1704896540
transform 1 0 74612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_702
timestamp 1704896540
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_714
timestamp 1704896540
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_726
timestamp 1704896540
transform 1 0 67804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_728
timestamp 1704896540
transform 1 0 67988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_740
timestamp 1704896540
transform 1 0 69092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_752
timestamp 1704896540
transform 1 0 70196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_764
timestamp 1704896540
transform 1 0 71300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_776
timestamp 1704896540
transform 1 0 72404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_782
timestamp 1704896540
transform 1 0 72956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_784
timestamp 1704896540
transform 1 0 73140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_796
timestamp 1704896540
transform 1 0 74244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_800
timestamp 1704896540
transform 1 0 74612 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_702
timestamp 1704896540
transform 1 0 65596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_714
timestamp 1704896540
transform 1 0 66700 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_726
timestamp 1704896540
transform 1 0 67804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_738
timestamp 1704896540
transform 1 0 68908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_750
timestamp 1704896540
transform 1 0 70012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_754
timestamp 1704896540
transform 1 0 70380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_756
timestamp 1704896540
transform 1 0 70564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_768
timestamp 1704896540
transform 1 0 71668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_780
timestamp 1704896540
transform 1 0 72772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_792
timestamp 1704896540
transform 1 0 73876 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_800
timestamp 1704896540
transform 1 0 74612 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_702
timestamp 1704896540
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_714
timestamp 1704896540
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_726
timestamp 1704896540
transform 1 0 67804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_728
timestamp 1704896540
transform 1 0 67988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_740
timestamp 1704896540
transform 1 0 69092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_752
timestamp 1704896540
transform 1 0 70196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_764
timestamp 1704896540
transform 1 0 71300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_776
timestamp 1704896540
transform 1 0 72404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_782
timestamp 1704896540
transform 1 0 72956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_784
timestamp 1704896540
transform 1 0 73140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_796
timestamp 1704896540
transform 1 0 74244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_800
timestamp 1704896540
transform 1 0 74612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_702
timestamp 1704896540
transform 1 0 65596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_714
timestamp 1704896540
transform 1 0 66700 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_726
timestamp 1704896540
transform 1 0 67804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_738
timestamp 1704896540
transform 1 0 68908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_750
timestamp 1704896540
transform 1 0 70012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_754
timestamp 1704896540
transform 1 0 70380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_756
timestamp 1704896540
transform 1 0 70564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_768
timestamp 1704896540
transform 1 0 71668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_780
timestamp 1704896540
transform 1 0 72772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_792
timestamp 1704896540
transform 1 0 73876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_800
timestamp 1704896540
transform 1 0 74612 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_702
timestamp 1704896540
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_714
timestamp 1704896540
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_726
timestamp 1704896540
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_728
timestamp 1704896540
transform 1 0 67988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_740
timestamp 1704896540
transform 1 0 69092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_752
timestamp 1704896540
transform 1 0 70196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_764
timestamp 1704896540
transform 1 0 71300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_776
timestamp 1704896540
transform 1 0 72404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_782
timestamp 1704896540
transform 1 0 72956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_784
timestamp 1704896540
transform 1 0 73140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_796
timestamp 1704896540
transform 1 0 74244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_800
timestamp 1704896540
transform 1 0 74612 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_702
timestamp 1704896540
transform 1 0 65596 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_714
timestamp 1704896540
transform 1 0 66700 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_726
timestamp 1704896540
transform 1 0 67804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_738
timestamp 1704896540
transform 1 0 68908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_750
timestamp 1704896540
transform 1 0 70012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_754
timestamp 1704896540
transform 1 0 70380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_756
timestamp 1704896540
transform 1 0 70564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_768
timestamp 1704896540
transform 1 0 71668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_780
timestamp 1704896540
transform 1 0 72772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_792
timestamp 1704896540
transform 1 0 73876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_800
timestamp 1704896540
transform 1 0 74612 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_702
timestamp 1704896540
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_714
timestamp 1704896540
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_726
timestamp 1704896540
transform 1 0 67804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_728
timestamp 1704896540
transform 1 0 67988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_740
timestamp 1704896540
transform 1 0 69092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_752
timestamp 1704896540
transform 1 0 70196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_764
timestamp 1704896540
transform 1 0 71300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_776
timestamp 1704896540
transform 1 0 72404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_782
timestamp 1704896540
transform 1 0 72956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_784
timestamp 1704896540
transform 1 0 73140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_796
timestamp 1704896540
transform 1 0 74244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_800
timestamp 1704896540
transform 1 0 74612 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_702
timestamp 1704896540
transform 1 0 65596 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_714
timestamp 1704896540
transform 1 0 66700 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_726
timestamp 1704896540
transform 1 0 67804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_738
timestamp 1704896540
transform 1 0 68908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_750
timestamp 1704896540
transform 1 0 70012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_754
timestamp 1704896540
transform 1 0 70380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_756
timestamp 1704896540
transform 1 0 70564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_768
timestamp 1704896540
transform 1 0 71668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_780
timestamp 1704896540
transform 1 0 72772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_792
timestamp 1704896540
transform 1 0 73876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_800
timestamp 1704896540
transform 1 0 74612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_702
timestamp 1704896540
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_714
timestamp 1704896540
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_726
timestamp 1704896540
transform 1 0 67804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_728
timestamp 1704896540
transform 1 0 67988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_740
timestamp 1704896540
transform 1 0 69092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_752
timestamp 1704896540
transform 1 0 70196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_764
timestamp 1704896540
transform 1 0 71300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_776
timestamp 1704896540
transform 1 0 72404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_782
timestamp 1704896540
transform 1 0 72956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_784
timestamp 1704896540
transform 1 0 73140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_796
timestamp 1704896540
transform 1 0 74244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_800
timestamp 1704896540
transform 1 0 74612 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_702
timestamp 1704896540
transform 1 0 65596 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_714
timestamp 1704896540
transform 1 0 66700 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_726
timestamp 1704896540
transform 1 0 67804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_738
timestamp 1704896540
transform 1 0 68908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_750
timestamp 1704896540
transform 1 0 70012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_754
timestamp 1704896540
transform 1 0 70380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_756
timestamp 1704896540
transform 1 0 70564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_768
timestamp 1704896540
transform 1 0 71668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_780
timestamp 1704896540
transform 1 0 72772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_792
timestamp 1704896540
transform 1 0 73876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_800
timestamp 1704896540
transform 1 0 74612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_702
timestamp 1704896540
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_714
timestamp 1704896540
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_726
timestamp 1704896540
transform 1 0 67804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_728
timestamp 1704896540
transform 1 0 67988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_740
timestamp 1704896540
transform 1 0 69092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_752
timestamp 1704896540
transform 1 0 70196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_764
timestamp 1704896540
transform 1 0 71300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_776
timestamp 1704896540
transform 1 0 72404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_782
timestamp 1704896540
transform 1 0 72956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_784
timestamp 1704896540
transform 1 0 73140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_796
timestamp 1704896540
transform 1 0 74244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_800
timestamp 1704896540
transform 1 0 74612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_702
timestamp 1704896540
transform 1 0 65596 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_714
timestamp 1704896540
transform 1 0 66700 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_726
timestamp 1704896540
transform 1 0 67804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_738
timestamp 1704896540
transform 1 0 68908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_750
timestamp 1704896540
transform 1 0 70012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_754
timestamp 1704896540
transform 1 0 70380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_756
timestamp 1704896540
transform 1 0 70564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_768
timestamp 1704896540
transform 1 0 71668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_780
timestamp 1704896540
transform 1 0 72772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_792
timestamp 1704896540
transform 1 0 73876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_800
timestamp 1704896540
transform 1 0 74612 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_702
timestamp 1704896540
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_714
timestamp 1704896540
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_726
timestamp 1704896540
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_728
timestamp 1704896540
transform 1 0 67988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_740
timestamp 1704896540
transform 1 0 69092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_752
timestamp 1704896540
transform 1 0 70196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_764
timestamp 1704896540
transform 1 0 71300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_776
timestamp 1704896540
transform 1 0 72404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_782
timestamp 1704896540
transform 1 0 72956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_784
timestamp 1704896540
transform 1 0 73140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_796
timestamp 1704896540
transform 1 0 74244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_800
timestamp 1704896540
transform 1 0 74612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_702
timestamp 1704896540
transform 1 0 65596 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_714
timestamp 1704896540
transform 1 0 66700 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_726
timestamp 1704896540
transform 1 0 67804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_738
timestamp 1704896540
transform 1 0 68908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_750
timestamp 1704896540
transform 1 0 70012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_754
timestamp 1704896540
transform 1 0 70380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_756
timestamp 1704896540
transform 1 0 70564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_768
timestamp 1704896540
transform 1 0 71668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_780
timestamp 1704896540
transform 1 0 72772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_792
timestamp 1704896540
transform 1 0 73876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_800
timestamp 1704896540
transform 1 0 74612 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_702
timestamp 1704896540
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_714
timestamp 1704896540
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_726
timestamp 1704896540
transform 1 0 67804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_728
timestamp 1704896540
transform 1 0 67988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_740
timestamp 1704896540
transform 1 0 69092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_752
timestamp 1704896540
transform 1 0 70196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_764
timestamp 1704896540
transform 1 0 71300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_776
timestamp 1704896540
transform 1 0 72404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_782
timestamp 1704896540
transform 1 0 72956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_784
timestamp 1704896540
transform 1 0 73140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_796
timestamp 1704896540
transform 1 0 74244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_800
timestamp 1704896540
transform 1 0 74612 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_702
timestamp 1704896540
transform 1 0 65596 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_714
timestamp 1704896540
transform 1 0 66700 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_726
timestamp 1704896540
transform 1 0 67804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_738
timestamp 1704896540
transform 1 0 68908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_750
timestamp 1704896540
transform 1 0 70012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_754
timestamp 1704896540
transform 1 0 70380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_756
timestamp 1704896540
transform 1 0 70564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_768
timestamp 1704896540
transform 1 0 71668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_780
timestamp 1704896540
transform 1 0 72772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_792
timestamp 1704896540
transform 1 0 73876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_800
timestamp 1704896540
transform 1 0 74612 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_702
timestamp 1704896540
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_714
timestamp 1704896540
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_726
timestamp 1704896540
transform 1 0 67804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_728
timestamp 1704896540
transform 1 0 67988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_740
timestamp 1704896540
transform 1 0 69092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_752
timestamp 1704896540
transform 1 0 70196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_764
timestamp 1704896540
transform 1 0 71300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_776
timestamp 1704896540
transform 1 0 72404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_782
timestamp 1704896540
transform 1 0 72956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_784
timestamp 1704896540
transform 1 0 73140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_796
timestamp 1704896540
transform 1 0 74244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_800
timestamp 1704896540
transform 1 0 74612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_702
timestamp 1704896540
transform 1 0 65596 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_714
timestamp 1704896540
transform 1 0 66700 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_726
timestamp 1704896540
transform 1 0 67804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_738
timestamp 1704896540
transform 1 0 68908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_750
timestamp 1704896540
transform 1 0 70012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_754
timestamp 1704896540
transform 1 0 70380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_756
timestamp 1704896540
transform 1 0 70564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_768
timestamp 1704896540
transform 1 0 71668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_780
timestamp 1704896540
transform 1 0 72772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_792
timestamp 1704896540
transform 1 0 73876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_800
timestamp 1704896540
transform 1 0 74612 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_702
timestamp 1704896540
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_714
timestamp 1704896540
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_726
timestamp 1704896540
transform 1 0 67804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_728
timestamp 1704896540
transform 1 0 67988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_740
timestamp 1704896540
transform 1 0 69092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_752
timestamp 1704896540
transform 1 0 70196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_764
timestamp 1704896540
transform 1 0 71300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_776
timestamp 1704896540
transform 1 0 72404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_782
timestamp 1704896540
transform 1 0 72956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_784
timestamp 1704896540
transform 1 0 73140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_796
timestamp 1704896540
transform 1 0 74244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_800
timestamp 1704896540
transform 1 0 74612 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_702
timestamp 1704896540
transform 1 0 65596 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_714
timestamp 1704896540
transform 1 0 66700 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_726
timestamp 1704896540
transform 1 0 67804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_738
timestamp 1704896540
transform 1 0 68908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_750
timestamp 1704896540
transform 1 0 70012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_754
timestamp 1704896540
transform 1 0 70380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_756
timestamp 1704896540
transform 1 0 70564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_768
timestamp 1704896540
transform 1 0 71668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_780
timestamp 1704896540
transform 1 0 72772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_792
timestamp 1704896540
transform 1 0 73876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_800
timestamp 1704896540
transform 1 0 74612 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_710
timestamp 1704896540
transform 1 0 66332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_722
timestamp 1704896540
transform 1 0 67436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_726
timestamp 1704896540
transform 1 0 67804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_728
timestamp 1704896540
transform 1 0 67988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_740
timestamp 1704896540
transform 1 0 69092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_752
timestamp 1704896540
transform 1 0 70196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_764
timestamp 1704896540
transform 1 0 71300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_776
timestamp 1704896540
transform 1 0 72404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_782
timestamp 1704896540
transform 1 0 72956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_784
timestamp 1704896540
transform 1 0 73140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_796
timestamp 1704896540
transform 1 0 74244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_800
timestamp 1704896540
transform 1 0 74612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_710
timestamp 1704896540
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_722
timestamp 1704896540
transform 1 0 67436 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_734
timestamp 1704896540
transform 1 0 68540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_746
timestamp 1704896540
transform 1 0 69644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_754
timestamp 1704896540
transform 1 0 70380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_756
timestamp 1704896540
transform 1 0 70564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_768
timestamp 1704896540
transform 1 0 71668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_780
timestamp 1704896540
transform 1 0 72772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_792
timestamp 1704896540
transform 1 0 73876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_800
timestamp 1704896540
transform 1 0 74612 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_710
timestamp 1704896540
transform 1 0 66332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_722
timestamp 1704896540
transform 1 0 67436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_726
timestamp 1704896540
transform 1 0 67804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_728
timestamp 1704896540
transform 1 0 67988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_740
timestamp 1704896540
transform 1 0 69092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_752
timestamp 1704896540
transform 1 0 70196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_764
timestamp 1704896540
transform 1 0 71300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_776
timestamp 1704896540
transform 1 0 72404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_782
timestamp 1704896540
transform 1 0 72956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_784
timestamp 1704896540
transform 1 0 73140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_796
timestamp 1704896540
transform 1 0 74244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_800
timestamp 1704896540
transform 1 0 74612 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_702
timestamp 1704896540
transform 1 0 65596 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_714
timestamp 1704896540
transform 1 0 66700 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_726
timestamp 1704896540
transform 1 0 67804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_738
timestamp 1704896540
transform 1 0 68908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_750
timestamp 1704896540
transform 1 0 70012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_754
timestamp 1704896540
transform 1 0 70380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_756
timestamp 1704896540
transform 1 0 70564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_768
timestamp 1704896540
transform 1 0 71668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_780
timestamp 1704896540
transform 1 0 72772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_792
timestamp 1704896540
transform 1 0 73876 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_800
timestamp 1704896540
transform 1 0 74612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_702
timestamp 1704896540
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_714
timestamp 1704896540
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_726
timestamp 1704896540
transform 1 0 67804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_728
timestamp 1704896540
transform 1 0 67988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_740
timestamp 1704896540
transform 1 0 69092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_752
timestamp 1704896540
transform 1 0 70196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_764
timestamp 1704896540
transform 1 0 71300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_776
timestamp 1704896540
transform 1 0 72404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_782
timestamp 1704896540
transform 1 0 72956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_784
timestamp 1704896540
transform 1 0 73140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_796
timestamp 1704896540
transform 1 0 74244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_800
timestamp 1704896540
transform 1 0 74612 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_702
timestamp 1704896540
transform 1 0 65596 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_714
timestamp 1704896540
transform 1 0 66700 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_726
timestamp 1704896540
transform 1 0 67804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_738
timestamp 1704896540
transform 1 0 68908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_750
timestamp 1704896540
transform 1 0 70012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_754
timestamp 1704896540
transform 1 0 70380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_756
timestamp 1704896540
transform 1 0 70564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_768
timestamp 1704896540
transform 1 0 71668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_780
timestamp 1704896540
transform 1 0 72772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_792
timestamp 1704896540
transform 1 0 73876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_800
timestamp 1704896540
transform 1 0 74612 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_710
timestamp 1704896540
transform 1 0 66332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_722
timestamp 1704896540
transform 1 0 67436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_726
timestamp 1704896540
transform 1 0 67804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_728
timestamp 1704896540
transform 1 0 67988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_740
timestamp 1704896540
transform 1 0 69092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_752
timestamp 1704896540
transform 1 0 70196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_764
timestamp 1704896540
transform 1 0 71300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_776
timestamp 1704896540
transform 1 0 72404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_782
timestamp 1704896540
transform 1 0 72956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_784
timestamp 1704896540
transform 1 0 73140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_796
timestamp 1704896540
transform 1 0 74244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_800
timestamp 1704896540
transform 1 0 74612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_718
timestamp 1704896540
transform 1 0 67068 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_730
timestamp 1704896540
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_742
timestamp 1704896540
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_754
timestamp 1704896540
transform 1 0 70380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_756
timestamp 1704896540
transform 1 0 70564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_768
timestamp 1704896540
transform 1 0 71668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_780
timestamp 1704896540
transform 1 0 72772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_792
timestamp 1704896540
transform 1 0 73876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_800
timestamp 1704896540
transform 1 0 74612 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_710
timestamp 1704896540
transform 1 0 66332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_722
timestamp 1704896540
transform 1 0 67436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_726
timestamp 1704896540
transform 1 0 67804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_728
timestamp 1704896540
transform 1 0 67988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_740
timestamp 1704896540
transform 1 0 69092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_752
timestamp 1704896540
transform 1 0 70196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_764
timestamp 1704896540
transform 1 0 71300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_776
timestamp 1704896540
transform 1 0 72404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_782
timestamp 1704896540
transform 1 0 72956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_784
timestamp 1704896540
transform 1 0 73140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_796
timestamp 1704896540
transform 1 0 74244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_800
timestamp 1704896540
transform 1 0 74612 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_702
timestamp 1704896540
transform 1 0 65596 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_714
timestamp 1704896540
transform 1 0 66700 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_726
timestamp 1704896540
transform 1 0 67804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_738
timestamp 1704896540
transform 1 0 68908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_750
timestamp 1704896540
transform 1 0 70012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_754
timestamp 1704896540
transform 1 0 70380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_756
timestamp 1704896540
transform 1 0 70564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_768
timestamp 1704896540
transform 1 0 71668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_780
timestamp 1704896540
transform 1 0 72772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_792
timestamp 1704896540
transform 1 0 73876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_800
timestamp 1704896540
transform 1 0 74612 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_710
timestamp 1704896540
transform 1 0 66332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_722
timestamp 1704896540
transform 1 0 67436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_726
timestamp 1704896540
transform 1 0 67804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_728
timestamp 1704896540
transform 1 0 67988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_740
timestamp 1704896540
transform 1 0 69092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_752
timestamp 1704896540
transform 1 0 70196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_764
timestamp 1704896540
transform 1 0 71300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_776
timestamp 1704896540
transform 1 0 72404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_782
timestamp 1704896540
transform 1 0 72956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_784
timestamp 1704896540
transform 1 0 73140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_796
timestamp 1704896540
transform 1 0 74244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_800
timestamp 1704896540
transform 1 0 74612 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_702
timestamp 1704896540
transform 1 0 65596 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_714
timestamp 1704896540
transform 1 0 66700 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_726
timestamp 1704896540
transform 1 0 67804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_738
timestamp 1704896540
transform 1 0 68908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_750
timestamp 1704896540
transform 1 0 70012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_754
timestamp 1704896540
transform 1 0 70380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_756
timestamp 1704896540
transform 1 0 70564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_768
timestamp 1704896540
transform 1 0 71668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_780
timestamp 1704896540
transform 1 0 72772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_792
timestamp 1704896540
transform 1 0 73876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_800
timestamp 1704896540
transform 1 0 74612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_710
timestamp 1704896540
transform 1 0 66332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_722
timestamp 1704896540
transform 1 0 67436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_726
timestamp 1704896540
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_728
timestamp 1704896540
transform 1 0 67988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_740
timestamp 1704896540
transform 1 0 69092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_752
timestamp 1704896540
transform 1 0 70196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_764
timestamp 1704896540
transform 1 0 71300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_776
timestamp 1704896540
transform 1 0 72404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_782
timestamp 1704896540
transform 1 0 72956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_784
timestamp 1704896540
transform 1 0 73140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_796
timestamp 1704896540
transform 1 0 74244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_800
timestamp 1704896540
transform 1 0 74612 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_702
timestamp 1704896540
transform 1 0 65596 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_714
timestamp 1704896540
transform 1 0 66700 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_726
timestamp 1704896540
transform 1 0 67804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_738
timestamp 1704896540
transform 1 0 68908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_750
timestamp 1704896540
transform 1 0 70012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_754
timestamp 1704896540
transform 1 0 70380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_756
timestamp 1704896540
transform 1 0 70564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_768
timestamp 1704896540
transform 1 0 71668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_780
timestamp 1704896540
transform 1 0 72772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_792
timestamp 1704896540
transform 1 0 73876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_800
timestamp 1704896540
transform 1 0 74612 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_710
timestamp 1704896540
transform 1 0 66332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_722
timestamp 1704896540
transform 1 0 67436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_726
timestamp 1704896540
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_728
timestamp 1704896540
transform 1 0 67988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_740
timestamp 1704896540
transform 1 0 69092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_752
timestamp 1704896540
transform 1 0 70196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_764
timestamp 1704896540
transform 1 0 71300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_776
timestamp 1704896540
transform 1 0 72404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_782
timestamp 1704896540
transform 1 0 72956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_784
timestamp 1704896540
transform 1 0 73140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_796
timestamp 1704896540
transform 1 0 74244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_800
timestamp 1704896540
transform 1 0 74612 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_702
timestamp 1704896540
transform 1 0 65596 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_714
timestamp 1704896540
transform 1 0 66700 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_726
timestamp 1704896540
transform 1 0 67804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_738
timestamp 1704896540
transform 1 0 68908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_750
timestamp 1704896540
transform 1 0 70012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_754
timestamp 1704896540
transform 1 0 70380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_756
timestamp 1704896540
transform 1 0 70564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_768
timestamp 1704896540
transform 1 0 71668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_780
timestamp 1704896540
transform 1 0 72772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_792
timestamp 1704896540
transform 1 0 73876 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_800
timestamp 1704896540
transform 1 0 74612 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_710
timestamp 1704896540
transform 1 0 66332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_722
timestamp 1704896540
transform 1 0 67436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_726
timestamp 1704896540
transform 1 0 67804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_728
timestamp 1704896540
transform 1 0 67988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_740
timestamp 1704896540
transform 1 0 69092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_752
timestamp 1704896540
transform 1 0 70196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_764
timestamp 1704896540
transform 1 0 71300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_776
timestamp 1704896540
transform 1 0 72404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_782
timestamp 1704896540
transform 1 0 72956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_784
timestamp 1704896540
transform 1 0 73140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_796
timestamp 1704896540
transform 1 0 74244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_800
timestamp 1704896540
transform 1 0 74612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_702
timestamp 1704896540
transform 1 0 65596 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_714
timestamp 1704896540
transform 1 0 66700 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_726
timestamp 1704896540
transform 1 0 67804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_738
timestamp 1704896540
transform 1 0 68908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_750
timestamp 1704896540
transform 1 0 70012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_754
timestamp 1704896540
transform 1 0 70380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_756
timestamp 1704896540
transform 1 0 70564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_768
timestamp 1704896540
transform 1 0 71668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_780
timestamp 1704896540
transform 1 0 72772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_792
timestamp 1704896540
transform 1 0 73876 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_800
timestamp 1704896540
transform 1 0 74612 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_710
timestamp 1704896540
transform 1 0 66332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_722
timestamp 1704896540
transform 1 0 67436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_726
timestamp 1704896540
transform 1 0 67804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_728
timestamp 1704896540
transform 1 0 67988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_740
timestamp 1704896540
transform 1 0 69092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_752
timestamp 1704896540
transform 1 0 70196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_764
timestamp 1704896540
transform 1 0 71300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_776
timestamp 1704896540
transform 1 0 72404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_782
timestamp 1704896540
transform 1 0 72956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_784
timestamp 1704896540
transform 1 0 73140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_796
timestamp 1704896540
transform 1 0 74244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_800
timestamp 1704896540
transform 1 0 74612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_710
timestamp 1704896540
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_722
timestamp 1704896540
transform 1 0 67436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_734
timestamp 1704896540
transform 1 0 68540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_746
timestamp 1704896540
transform 1 0 69644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_754
timestamp 1704896540
transform 1 0 70380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_756
timestamp 1704896540
transform 1 0 70564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_768
timestamp 1704896540
transform 1 0 71668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_780
timestamp 1704896540
transform 1 0 72772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_792
timestamp 1704896540
transform 1 0 73876 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_800
timestamp 1704896540
transform 1 0 74612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_722
timestamp 1704896540
transform 1 0 67436 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_726
timestamp 1704896540
transform 1 0 67804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_728
timestamp 1704896540
transform 1 0 67988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_740
timestamp 1704896540
transform 1 0 69092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_752
timestamp 1704896540
transform 1 0 70196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_764
timestamp 1704896540
transform 1 0 71300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_776
timestamp 1704896540
transform 1 0 72404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_782
timestamp 1704896540
transform 1 0 72956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_784
timestamp 1704896540
transform 1 0 73140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_796
timestamp 1704896540
transform 1 0 74244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_800
timestamp 1704896540
transform 1 0 74612 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_702
timestamp 1704896540
transform 1 0 65596 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_714
timestamp 1704896540
transform 1 0 66700 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_726
timestamp 1704896540
transform 1 0 67804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_738
timestamp 1704896540
transform 1 0 68908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_750
timestamp 1704896540
transform 1 0 70012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_754
timestamp 1704896540
transform 1 0 70380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_756
timestamp 1704896540
transform 1 0 70564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_768
timestamp 1704896540
transform 1 0 71668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_780
timestamp 1704896540
transform 1 0 72772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_792
timestamp 1704896540
transform 1 0 73876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_800
timestamp 1704896540
transform 1 0 74612 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_710
timestamp 1704896540
transform 1 0 66332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_722
timestamp 1704896540
transform 1 0 67436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_726
timestamp 1704896540
transform 1 0 67804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_728
timestamp 1704896540
transform 1 0 67988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_740
timestamp 1704896540
transform 1 0 69092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_752
timestamp 1704896540
transform 1 0 70196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_764
timestamp 1704896540
transform 1 0 71300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_776
timestamp 1704896540
transform 1 0 72404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_782
timestamp 1704896540
transform 1 0 72956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_784
timestamp 1704896540
transform 1 0 73140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_796
timestamp 1704896540
transform 1 0 74244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_800
timestamp 1704896540
transform 1 0 74612 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_718
timestamp 1704896540
transform 1 0 67068 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_730
timestamp 1704896540
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_742
timestamp 1704896540
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_754
timestamp 1704896540
transform 1 0 70380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_756
timestamp 1704896540
transform 1 0 70564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_768
timestamp 1704896540
transform 1 0 71668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_780
timestamp 1704896540
transform 1 0 72772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_792
timestamp 1704896540
transform 1 0 73876 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_800
timestamp 1704896540
transform 1 0 74612 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_710
timestamp 1704896540
transform 1 0 66332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_722
timestamp 1704896540
transform 1 0 67436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_726
timestamp 1704896540
transform 1 0 67804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_728
timestamp 1704896540
transform 1 0 67988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_740
timestamp 1704896540
transform 1 0 69092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_752
timestamp 1704896540
transform 1 0 70196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_764
timestamp 1704896540
transform 1 0 71300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_776
timestamp 1704896540
transform 1 0 72404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_782
timestamp 1704896540
transform 1 0 72956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_784
timestamp 1704896540
transform 1 0 73140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_796
timestamp 1704896540
transform 1 0 74244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_800
timestamp 1704896540
transform 1 0 74612 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_702
timestamp 1704896540
transform 1 0 65596 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_714
timestamp 1704896540
transform 1 0 66700 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_726
timestamp 1704896540
transform 1 0 67804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_738
timestamp 1704896540
transform 1 0 68908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_750
timestamp 1704896540
transform 1 0 70012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_754
timestamp 1704896540
transform 1 0 70380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_756
timestamp 1704896540
transform 1 0 70564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_768
timestamp 1704896540
transform 1 0 71668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_780
timestamp 1704896540
transform 1 0 72772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_792
timestamp 1704896540
transform 1 0 73876 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_800
timestamp 1704896540
transform 1 0 74612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_710
timestamp 1704896540
transform 1 0 66332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_722
timestamp 1704896540
transform 1 0 67436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_726
timestamp 1704896540
transform 1 0 67804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_728
timestamp 1704896540
transform 1 0 67988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_740
timestamp 1704896540
transform 1 0 69092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_752
timestamp 1704896540
transform 1 0 70196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_764
timestamp 1704896540
transform 1 0 71300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_776
timestamp 1704896540
transform 1 0 72404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_782
timestamp 1704896540
transform 1 0 72956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_784
timestamp 1704896540
transform 1 0 73140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_796
timestamp 1704896540
transform 1 0 74244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_800
timestamp 1704896540
transform 1 0 74612 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_702
timestamp 1704896540
transform 1 0 65596 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_714
timestamp 1704896540
transform 1 0 66700 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_726
timestamp 1704896540
transform 1 0 67804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_738
timestamp 1704896540
transform 1 0 68908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_750
timestamp 1704896540
transform 1 0 70012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_754
timestamp 1704896540
transform 1 0 70380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_756
timestamp 1704896540
transform 1 0 70564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_768
timestamp 1704896540
transform 1 0 71668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_780
timestamp 1704896540
transform 1 0 72772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_792
timestamp 1704896540
transform 1 0 73876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_800
timestamp 1704896540
transform 1 0 74612 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_710
timestamp 1704896540
transform 1 0 66332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_722
timestamp 1704896540
transform 1 0 67436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_726
timestamp 1704896540
transform 1 0 67804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_728
timestamp 1704896540
transform 1 0 67988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_740
timestamp 1704896540
transform 1 0 69092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_752
timestamp 1704896540
transform 1 0 70196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_764
timestamp 1704896540
transform 1 0 71300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_776
timestamp 1704896540
transform 1 0 72404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_782
timestamp 1704896540
transform 1 0 72956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_784
timestamp 1704896540
transform 1 0 73140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_796
timestamp 1704896540
transform 1 0 74244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_800
timestamp 1704896540
transform 1 0 74612 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_702
timestamp 1704896540
transform 1 0 65596 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_714
timestamp 1704896540
transform 1 0 66700 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_726
timestamp 1704896540
transform 1 0 67804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_738
timestamp 1704896540
transform 1 0 68908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_750
timestamp 1704896540
transform 1 0 70012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_754
timestamp 1704896540
transform 1 0 70380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_756
timestamp 1704896540
transform 1 0 70564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_768
timestamp 1704896540
transform 1 0 71668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_780
timestamp 1704896540
transform 1 0 72772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_792
timestamp 1704896540
transform 1 0 73876 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_800
timestamp 1704896540
transform 1 0 74612 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_710
timestamp 1704896540
transform 1 0 66332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_722
timestamp 1704896540
transform 1 0 67436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_726
timestamp 1704896540
transform 1 0 67804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_728
timestamp 1704896540
transform 1 0 67988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_740
timestamp 1704896540
transform 1 0 69092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_752
timestamp 1704896540
transform 1 0 70196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_764
timestamp 1704896540
transform 1 0 71300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_776
timestamp 1704896540
transform 1 0 72404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_782
timestamp 1704896540
transform 1 0 72956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_784
timestamp 1704896540
transform 1 0 73140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_796
timestamp 1704896540
transform 1 0 74244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_800
timestamp 1704896540
transform 1 0 74612 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_702
timestamp 1704896540
transform 1 0 65596 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_714
timestamp 1704896540
transform 1 0 66700 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_726
timestamp 1704896540
transform 1 0 67804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_738
timestamp 1704896540
transform 1 0 68908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_750
timestamp 1704896540
transform 1 0 70012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_754
timestamp 1704896540
transform 1 0 70380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_756
timestamp 1704896540
transform 1 0 70564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_768
timestamp 1704896540
transform 1 0 71668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_780
timestamp 1704896540
transform 1 0 72772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_792
timestamp 1704896540
transform 1 0 73876 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_800
timestamp 1704896540
transform 1 0 74612 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_702
timestamp 1704896540
transform 1 0 65596 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_710
timestamp 1704896540
transform 1 0 66332 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_719
timestamp 1704896540
transform 1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_728
timestamp 1704896540
transform 1 0 67988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_740
timestamp 1704896540
transform 1 0 69092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_752
timestamp 1704896540
transform 1 0 70196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_764
timestamp 1704896540
transform 1 0 71300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_776
timestamp 1704896540
transform 1 0 72404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_782
timestamp 1704896540
transform 1 0 72956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_784
timestamp 1704896540
transform 1 0 73140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_796
timestamp 1704896540
transform 1 0 74244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_800
timestamp 1704896540
transform 1 0 74612 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_702
timestamp 1704896540
transform 1 0 65596 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_714
timestamp 1704896540
transform 1 0 66700 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_726
timestamp 1704896540
transform 1 0 67804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_738
timestamp 1704896540
transform 1 0 68908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_750
timestamp 1704896540
transform 1 0 70012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_754
timestamp 1704896540
transform 1 0 70380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_756
timestamp 1704896540
transform 1 0 70564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_768
timestamp 1704896540
transform 1 0 71668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_780
timestamp 1704896540
transform 1 0 72772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_792
timestamp 1704896540
transform 1 0 73876 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_800
timestamp 1704896540
transform 1 0 74612 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_702
timestamp 1704896540
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_714
timestamp 1704896540
transform 1 0 66700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_726
timestamp 1704896540
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_728
timestamp 1704896540
transform 1 0 67988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_740
timestamp 1704896540
transform 1 0 69092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_752
timestamp 1704896540
transform 1 0 70196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_764
timestamp 1704896540
transform 1 0 71300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_776
timestamp 1704896540
transform 1 0 72404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_782
timestamp 1704896540
transform 1 0 72956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_784
timestamp 1704896540
transform 1 0 73140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_796
timestamp 1704896540
transform 1 0 74244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_800
timestamp 1704896540
transform 1 0 74612 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_702
timestamp 1704896540
transform 1 0 65596 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_714
timestamp 1704896540
transform 1 0 66700 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_726
timestamp 1704896540
transform 1 0 67804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_738
timestamp 1704896540
transform 1 0 68908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_750
timestamp 1704896540
transform 1 0 70012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_754
timestamp 1704896540
transform 1 0 70380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_756
timestamp 1704896540
transform 1 0 70564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_768
timestamp 1704896540
transform 1 0 71668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_780
timestamp 1704896540
transform 1 0 72772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_792
timestamp 1704896540
transform 1 0 73876 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_800
timestamp 1704896540
transform 1 0 74612 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_705
timestamp 1704896540
transform 1 0 65872 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_717
timestamp 1704896540
transform 1 0 66976 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_725
timestamp 1704896540
transform 1 0 67712 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_736
timestamp 1704896540
transform 1 0 68724 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_748
timestamp 1704896540
transform 1 0 69828 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_760
timestamp 1704896540
transform 1 0 70932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_772
timestamp 1704896540
transform 1 0 72036 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_780
timestamp 1704896540
transform 1 0 72772 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_784
timestamp 1704896540
transform 1 0 73140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_796
timestamp 1704896540
transform 1 0 74244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_800
timestamp 1704896540
transform 1 0 74612 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_702
timestamp 1704896540
transform 1 0 65596 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_714
timestamp 1704896540
transform 1 0 66700 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_726
timestamp 1704896540
transform 1 0 67804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_738
timestamp 1704896540
transform 1 0 68908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_750
timestamp 1704896540
transform 1 0 70012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_754
timestamp 1704896540
transform 1 0 70380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_756
timestamp 1704896540
transform 1 0 70564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_768
timestamp 1704896540
transform 1 0 71668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_780
timestamp 1704896540
transform 1 0 72772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_792
timestamp 1704896540
transform 1 0 73876 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_800
timestamp 1704896540
transform 1 0 74612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_705
timestamp 1704896540
transform 1 0 65872 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_717
timestamp 1704896540
transform 1 0 66976 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_725
timestamp 1704896540
transform 1 0 67712 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_728
timestamp 1704896540
transform 1 0 67988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_740
timestamp 1704896540
transform 1 0 69092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_752
timestamp 1704896540
transform 1 0 70196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_764
timestamp 1704896540
transform 1 0 71300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_776
timestamp 1704896540
transform 1 0 72404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_782
timestamp 1704896540
transform 1 0 72956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_784
timestamp 1704896540
transform 1 0 73140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_796
timestamp 1704896540
transform 1 0 74244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_800
timestamp 1704896540
transform 1 0 74612 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_702
timestamp 1704896540
transform 1 0 65596 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_714
timestamp 1704896540
transform 1 0 66700 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_726
timestamp 1704896540
transform 1 0 67804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_738
timestamp 1704896540
transform 1 0 68908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_750
timestamp 1704896540
transform 1 0 70012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_754
timestamp 1704896540
transform 1 0 70380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_756
timestamp 1704896540
transform 1 0 70564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_768
timestamp 1704896540
transform 1 0 71668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_780
timestamp 1704896540
transform 1 0 72772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_792
timestamp 1704896540
transform 1 0 73876 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_800
timestamp 1704896540
transform 1 0 74612 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_702
timestamp 1704896540
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_714
timestamp 1704896540
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_726
timestamp 1704896540
transform 1 0 67804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_728
timestamp 1704896540
transform 1 0 67988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_740
timestamp 1704896540
transform 1 0 69092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_752
timestamp 1704896540
transform 1 0 70196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_764
timestamp 1704896540
transform 1 0 71300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_776
timestamp 1704896540
transform 1 0 72404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_782
timestamp 1704896540
transform 1 0 72956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_784
timestamp 1704896540
transform 1 0 73140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_796
timestamp 1704896540
transform 1 0 74244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_800
timestamp 1704896540
transform 1 0 74612 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_702
timestamp 1704896540
transform 1 0 65596 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_714
timestamp 1704896540
transform 1 0 66700 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_726
timestamp 1704896540
transform 1 0 67804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_738
timestamp 1704896540
transform 1 0 68908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_750
timestamp 1704896540
transform 1 0 70012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_754
timestamp 1704896540
transform 1 0 70380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_756
timestamp 1704896540
transform 1 0 70564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_768
timestamp 1704896540
transform 1 0 71668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_780
timestamp 1704896540
transform 1 0 72772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_792
timestamp 1704896540
transform 1 0 73876 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_800
timestamp 1704896540
transform 1 0 74612 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_702
timestamp 1704896540
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_714
timestamp 1704896540
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_726
timestamp 1704896540
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_728
timestamp 1704896540
transform 1 0 67988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_740
timestamp 1704896540
transform 1 0 69092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_752
timestamp 1704896540
transform 1 0 70196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_764
timestamp 1704896540
transform 1 0 71300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_776
timestamp 1704896540
transform 1 0 72404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_782
timestamp 1704896540
transform 1 0 72956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_784
timestamp 1704896540
transform 1 0 73140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_796
timestamp 1704896540
transform 1 0 74244 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_800
timestamp 1704896540
transform 1 0 74612 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_702
timestamp 1704896540
transform 1 0 65596 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_714
timestamp 1704896540
transform 1 0 66700 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_726
timestamp 1704896540
transform 1 0 67804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_738
timestamp 1704896540
transform 1 0 68908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_750
timestamp 1704896540
transform 1 0 70012 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_754
timestamp 1704896540
transform 1 0 70380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_756
timestamp 1704896540
transform 1 0 70564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_768
timestamp 1704896540
transform 1 0 71668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_780
timestamp 1704896540
transform 1 0 72772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_792
timestamp 1704896540
transform 1 0 73876 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_800
timestamp 1704896540
transform 1 0 74612 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_708
timestamp 1704896540
transform 1 0 66148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_720
timestamp 1704896540
transform 1 0 67252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_726
timestamp 1704896540
transform 1 0 67804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_728
timestamp 1704896540
transform 1 0 67988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_740
timestamp 1704896540
transform 1 0 69092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_752
timestamp 1704896540
transform 1 0 70196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_764
timestamp 1704896540
transform 1 0 71300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_776
timestamp 1704896540
transform 1 0 72404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_782
timestamp 1704896540
transform 1 0 72956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_784
timestamp 1704896540
transform 1 0 73140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_84_796
timestamp 1704896540
transform 1 0 74244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_800
timestamp 1704896540
transform 1 0 74612 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_702
timestamp 1704896540
transform 1 0 65596 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_714
timestamp 1704896540
transform 1 0 66700 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_726
timestamp 1704896540
transform 1 0 67804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_738
timestamp 1704896540
transform 1 0 68908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_750
timestamp 1704896540
transform 1 0 70012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_754
timestamp 1704896540
transform 1 0 70380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_756
timestamp 1704896540
transform 1 0 70564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_768
timestamp 1704896540
transform 1 0 71668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_780
timestamp 1704896540
transform 1 0 72772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_792
timestamp 1704896540
transform 1 0 73876 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_800
timestamp 1704896540
transform 1 0 74612 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_702
timestamp 1704896540
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_714
timestamp 1704896540
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_726
timestamp 1704896540
transform 1 0 67804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_728
timestamp 1704896540
transform 1 0 67988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_740
timestamp 1704896540
transform 1 0 69092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_752
timestamp 1704896540
transform 1 0 70196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_764
timestamp 1704896540
transform 1 0 71300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_776
timestamp 1704896540
transform 1 0 72404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_782
timestamp 1704896540
transform 1 0 72956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_784
timestamp 1704896540
transform 1 0 73140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86_796
timestamp 1704896540
transform 1 0 74244 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_800
timestamp 1704896540
transform 1 0 74612 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_702
timestamp 1704896540
transform 1 0 65596 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_714
timestamp 1704896540
transform 1 0 66700 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_726
timestamp 1704896540
transform 1 0 67804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_738
timestamp 1704896540
transform 1 0 68908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_750
timestamp 1704896540
transform 1 0 70012 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_754
timestamp 1704896540
transform 1 0 70380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_756
timestamp 1704896540
transform 1 0 70564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_768
timestamp 1704896540
transform 1 0 71668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_780
timestamp 1704896540
transform 1 0 72772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_792
timestamp 1704896540
transform 1 0 73876 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_800
timestamp 1704896540
transform 1 0 74612 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_705
timestamp 1704896540
transform 1 0 65872 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_717
timestamp 1704896540
transform 1 0 66976 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88_725
timestamp 1704896540
transform 1 0 67712 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_728
timestamp 1704896540
transform 1 0 67988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_740
timestamp 1704896540
transform 1 0 69092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_752
timestamp 1704896540
transform 1 0 70196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_764
timestamp 1704896540
transform 1 0 71300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_776
timestamp 1704896540
transform 1 0 72404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_782
timestamp 1704896540
transform 1 0 72956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_784
timestamp 1704896540
transform 1 0 73140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88_796
timestamp 1704896540
transform 1 0 74244 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_800
timestamp 1704896540
transform 1 0 74612 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_705
timestamp 1704896540
transform 1 0 65872 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_717
timestamp 1704896540
transform 1 0 66976 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_729
timestamp 1704896540
transform 1 0 68080 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_741
timestamp 1704896540
transform 1 0 69184 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_753
timestamp 1704896540
transform 1 0 70288 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_756
timestamp 1704896540
transform 1 0 70564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_768
timestamp 1704896540
transform 1 0 71668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_780
timestamp 1704896540
transform 1 0 72772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_792
timestamp 1704896540
transform 1 0 73876 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_800
timestamp 1704896540
transform 1 0 74612 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_705
timestamp 1704896540
transform 1 0 65872 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_717
timestamp 1704896540
transform 1 0 66976 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_725
timestamp 1704896540
transform 1 0 67712 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_728
timestamp 1704896540
transform 1 0 67988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_740
timestamp 1704896540
transform 1 0 69092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_752
timestamp 1704896540
transform 1 0 70196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_764
timestamp 1704896540
transform 1 0 71300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_776
timestamp 1704896540
transform 1 0 72404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_782
timestamp 1704896540
transform 1 0 72956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_784
timestamp 1704896540
transform 1 0 73140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90_796
timestamp 1704896540
transform 1 0 74244 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_800
timestamp 1704896540
transform 1 0 74612 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_702
timestamp 1704896540
transform 1 0 65596 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_714
timestamp 1704896540
transform 1 0 66700 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_726
timestamp 1704896540
transform 1 0 67804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_738
timestamp 1704896540
transform 1 0 68908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_750
timestamp 1704896540
transform 1 0 70012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_754
timestamp 1704896540
transform 1 0 70380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_756
timestamp 1704896540
transform 1 0 70564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_768
timestamp 1704896540
transform 1 0 71668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_780
timestamp 1704896540
transform 1 0 72772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_792
timestamp 1704896540
transform 1 0 73876 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_800
timestamp 1704896540
transform 1 0 74612 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_702
timestamp 1704896540
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_714
timestamp 1704896540
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_726
timestamp 1704896540
transform 1 0 67804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_728
timestamp 1704896540
transform 1 0 67988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_740
timestamp 1704896540
transform 1 0 69092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_752
timestamp 1704896540
transform 1 0 70196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_764
timestamp 1704896540
transform 1 0 71300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_776
timestamp 1704896540
transform 1 0 72404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_782
timestamp 1704896540
transform 1 0 72956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_784
timestamp 1704896540
transform 1 0 73140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92_796
timestamp 1704896540
transform 1 0 74244 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_800
timestamp 1704896540
transform 1 0 74612 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_702
timestamp 1704896540
transform 1 0 65596 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_714
timestamp 1704896540
transform 1 0 66700 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_726
timestamp 1704896540
transform 1 0 67804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_738
timestamp 1704896540
transform 1 0 68908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_750
timestamp 1704896540
transform 1 0 70012 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_754
timestamp 1704896540
transform 1 0 70380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_756
timestamp 1704896540
transform 1 0 70564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_768
timestamp 1704896540
transform 1 0 71668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_780
timestamp 1704896540
transform 1 0 72772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_792
timestamp 1704896540
transform 1 0 73876 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_800
timestamp 1704896540
transform 1 0 74612 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_708
timestamp 1704896540
transform 1 0 66148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_720
timestamp 1704896540
transform 1 0 67252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_726
timestamp 1704896540
transform 1 0 67804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_728
timestamp 1704896540
transform 1 0 67988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_740
timestamp 1704896540
transform 1 0 69092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_752
timestamp 1704896540
transform 1 0 70196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_764
timestamp 1704896540
transform 1 0 71300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_776
timestamp 1704896540
transform 1 0 72404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_782
timestamp 1704896540
transform 1 0 72956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_784
timestamp 1704896540
transform 1 0 73140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_796
timestamp 1704896540
transform 1 0 74244 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_800
timestamp 1704896540
transform 1 0 74612 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_702
timestamp 1704896540
transform 1 0 65596 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_714
timestamp 1704896540
transform 1 0 66700 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_726
timestamp 1704896540
transform 1 0 67804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_738
timestamp 1704896540
transform 1 0 68908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_750
timestamp 1704896540
transform 1 0 70012 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_754
timestamp 1704896540
transform 1 0 70380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_756
timestamp 1704896540
transform 1 0 70564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_768
timestamp 1704896540
transform 1 0 71668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_780
timestamp 1704896540
transform 1 0 72772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_792
timestamp 1704896540
transform 1 0 73876 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_800
timestamp 1704896540
transform 1 0 74612 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_702
timestamp 1704896540
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_714
timestamp 1704896540
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_726
timestamp 1704896540
transform 1 0 67804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_728
timestamp 1704896540
transform 1 0 67988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_740
timestamp 1704896540
transform 1 0 69092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_752
timestamp 1704896540
transform 1 0 70196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_764
timestamp 1704896540
transform 1 0 71300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_776
timestamp 1704896540
transform 1 0 72404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_782
timestamp 1704896540
transform 1 0 72956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_784
timestamp 1704896540
transform 1 0 73140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_796
timestamp 1704896540
transform 1 0 74244 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_800
timestamp 1704896540
transform 1 0 74612 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_702
timestamp 1704896540
transform 1 0 65596 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_714
timestamp 1704896540
transform 1 0 66700 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_726
timestamp 1704896540
transform 1 0 67804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_738
timestamp 1704896540
transform 1 0 68908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_750
timestamp 1704896540
transform 1 0 70012 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_754
timestamp 1704896540
transform 1 0 70380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_756
timestamp 1704896540
transform 1 0 70564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_768
timestamp 1704896540
transform 1 0 71668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_780
timestamp 1704896540
transform 1 0 72772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_792
timestamp 1704896540
transform 1 0 73876 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_800
timestamp 1704896540
transform 1 0 74612 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_702
timestamp 1704896540
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_714
timestamp 1704896540
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_726
timestamp 1704896540
transform 1 0 67804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_728
timestamp 1704896540
transform 1 0 67988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_740
timestamp 1704896540
transform 1 0 69092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_752
timestamp 1704896540
transform 1 0 70196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_764
timestamp 1704896540
transform 1 0 71300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_776
timestamp 1704896540
transform 1 0 72404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_782
timestamp 1704896540
transform 1 0 72956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_784
timestamp 1704896540
transform 1 0 73140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_796
timestamp 1704896540
transform 1 0 74244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_800
timestamp 1704896540
transform 1 0 74612 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_702
timestamp 1704896540
transform 1 0 65596 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_714
timestamp 1704896540
transform 1 0 66700 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_726
timestamp 1704896540
transform 1 0 67804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_738
timestamp 1704896540
transform 1 0 68908 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_750
timestamp 1704896540
transform 1 0 70012 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_754
timestamp 1704896540
transform 1 0 70380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_756
timestamp 1704896540
transform 1 0 70564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_768
timestamp 1704896540
transform 1 0 71668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_780
timestamp 1704896540
transform 1 0 72772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_792
timestamp 1704896540
transform 1 0 73876 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_800
timestamp 1704896540
transform 1 0 74612 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_702
timestamp 1704896540
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_714
timestamp 1704896540
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_726
timestamp 1704896540
transform 1 0 67804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_728
timestamp 1704896540
transform 1 0 67988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_740
timestamp 1704896540
transform 1 0 69092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_752
timestamp 1704896540
transform 1 0 70196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_764
timestamp 1704896540
transform 1 0 71300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_776
timestamp 1704896540
transform 1 0 72404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_782
timestamp 1704896540
transform 1 0 72956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_784
timestamp 1704896540
transform 1 0 73140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_796
timestamp 1704896540
transform 1 0 74244 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_800
timestamp 1704896540
transform 1 0 74612 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_702
timestamp 1704896540
transform 1 0 65596 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_714
timestamp 1704896540
transform 1 0 66700 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_726
timestamp 1704896540
transform 1 0 67804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_738
timestamp 1704896540
transform 1 0 68908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_750
timestamp 1704896540
transform 1 0 70012 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_754
timestamp 1704896540
transform 1 0 70380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_756
timestamp 1704896540
transform 1 0 70564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_768
timestamp 1704896540
transform 1 0 71668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_780
timestamp 1704896540
transform 1 0 72772 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_792
timestamp 1704896540
transform 1 0 73876 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_800
timestamp 1704896540
transform 1 0 74612 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_702
timestamp 1704896540
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_714
timestamp 1704896540
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_726
timestamp 1704896540
transform 1 0 67804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_728
timestamp 1704896540
transform 1 0 67988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_740
timestamp 1704896540
transform 1 0 69092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_752
timestamp 1704896540
transform 1 0 70196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_764
timestamp 1704896540
transform 1 0 71300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_776
timestamp 1704896540
transform 1 0 72404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_782
timestamp 1704896540
transform 1 0 72956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_784
timestamp 1704896540
transform 1 0 73140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_796
timestamp 1704896540
transform 1 0 74244 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_800
timestamp 1704896540
transform 1 0 74612 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_702
timestamp 1704896540
transform 1 0 65596 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_714
timestamp 1704896540
transform 1 0 66700 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_726
timestamp 1704896540
transform 1 0 67804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_738
timestamp 1704896540
transform 1 0 68908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_750
timestamp 1704896540
transform 1 0 70012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_754
timestamp 1704896540
transform 1 0 70380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_756
timestamp 1704896540
transform 1 0 70564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_768
timestamp 1704896540
transform 1 0 71668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_780
timestamp 1704896540
transform 1 0 72772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_792
timestamp 1704896540
transform 1 0 73876 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_800
timestamp 1704896540
transform 1 0 74612 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_702
timestamp 1704896540
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_714
timestamp 1704896540
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_726
timestamp 1704896540
transform 1 0 67804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_728
timestamp 1704896540
transform 1 0 67988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_740
timestamp 1704896540
transform 1 0 69092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_752
timestamp 1704896540
transform 1 0 70196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_764
timestamp 1704896540
transform 1 0 71300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_776
timestamp 1704896540
transform 1 0 72404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_782
timestamp 1704896540
transform 1 0 72956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_784
timestamp 1704896540
transform 1 0 73140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_796
timestamp 1704896540
transform 1 0 74244 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_800
timestamp 1704896540
transform 1 0 74612 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_702
timestamp 1704896540
transform 1 0 65596 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_714
timestamp 1704896540
transform 1 0 66700 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_726
timestamp 1704896540
transform 1 0 67804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_738
timestamp 1704896540
transform 1 0 68908 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_750
timestamp 1704896540
transform 1 0 70012 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_754
timestamp 1704896540
transform 1 0 70380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_756
timestamp 1704896540
transform 1 0 70564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_768
timestamp 1704896540
transform 1 0 71668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_780
timestamp 1704896540
transform 1 0 72772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_792
timestamp 1704896540
transform 1 0 73876 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_800
timestamp 1704896540
transform 1 0 74612 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_702
timestamp 1704896540
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_714
timestamp 1704896540
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_726
timestamp 1704896540
transform 1 0 67804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_728
timestamp 1704896540
transform 1 0 67988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_740
timestamp 1704896540
transform 1 0 69092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_752
timestamp 1704896540
transform 1 0 70196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_764
timestamp 1704896540
transform 1 0 71300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_776
timestamp 1704896540
transform 1 0 72404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_782
timestamp 1704896540
transform 1 0 72956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_784
timestamp 1704896540
transform 1 0 73140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106_796
timestamp 1704896540
transform 1 0 74244 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_800
timestamp 1704896540
transform 1 0 74612 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_702
timestamp 1704896540
transform 1 0 65596 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_714
timestamp 1704896540
transform 1 0 66700 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_726
timestamp 1704896540
transform 1 0 67804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_738
timestamp 1704896540
transform 1 0 68908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_750
timestamp 1704896540
transform 1 0 70012 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_754
timestamp 1704896540
transform 1 0 70380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_756
timestamp 1704896540
transform 1 0 70564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_768
timestamp 1704896540
transform 1 0 71668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_780
timestamp 1704896540
transform 1 0 72772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_792
timestamp 1704896540
transform 1 0 73876 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_800
timestamp 1704896540
transform 1 0 74612 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_702
timestamp 1704896540
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_714
timestamp 1704896540
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_726
timestamp 1704896540
transform 1 0 67804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_728
timestamp 1704896540
transform 1 0 67988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_740
timestamp 1704896540
transform 1 0 69092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_752
timestamp 1704896540
transform 1 0 70196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_764
timestamp 1704896540
transform 1 0 71300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_776
timestamp 1704896540
transform 1 0 72404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_782
timestamp 1704896540
transform 1 0 72956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_784
timestamp 1704896540
transform 1 0 73140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108_796
timestamp 1704896540
transform 1 0 74244 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_800
timestamp 1704896540
transform 1 0 74612 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_702
timestamp 1704896540
transform 1 0 65596 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_714
timestamp 1704896540
transform 1 0 66700 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_726
timestamp 1704896540
transform 1 0 67804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_738
timestamp 1704896540
transform 1 0 68908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_750
timestamp 1704896540
transform 1 0 70012 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_754
timestamp 1704896540
transform 1 0 70380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_756
timestamp 1704896540
transform 1 0 70564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_768
timestamp 1704896540
transform 1 0 71668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_780
timestamp 1704896540
transform 1 0 72772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_792
timestamp 1704896540
transform 1 0 73876 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_800
timestamp 1704896540
transform 1 0 74612 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_702
timestamp 1704896540
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_714
timestamp 1704896540
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_726
timestamp 1704896540
transform 1 0 67804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_728
timestamp 1704896540
transform 1 0 67988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_740
timestamp 1704896540
transform 1 0 69092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_752
timestamp 1704896540
transform 1 0 70196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_764
timestamp 1704896540
transform 1 0 71300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_776
timestamp 1704896540
transform 1 0 72404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_782
timestamp 1704896540
transform 1 0 72956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_784
timestamp 1704896540
transform 1 0 73140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_796
timestamp 1704896540
transform 1 0 74244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_800
timestamp 1704896540
transform 1 0 74612 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_702
timestamp 1704896540
transform 1 0 65596 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_714
timestamp 1704896540
transform 1 0 66700 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_726
timestamp 1704896540
transform 1 0 67804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_738
timestamp 1704896540
transform 1 0 68908 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_750
timestamp 1704896540
transform 1 0 70012 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_754
timestamp 1704896540
transform 1 0 70380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_756
timestamp 1704896540
transform 1 0 70564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_768
timestamp 1704896540
transform 1 0 71668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_780
timestamp 1704896540
transform 1 0 72772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_792
timestamp 1704896540
transform 1 0 73876 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_800
timestamp 1704896540
transform 1 0 74612 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_702
timestamp 1704896540
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_714
timestamp 1704896540
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_726
timestamp 1704896540
transform 1 0 67804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_728
timestamp 1704896540
transform 1 0 67988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_740
timestamp 1704896540
transform 1 0 69092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_752
timestamp 1704896540
transform 1 0 70196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_764
timestamp 1704896540
transform 1 0 71300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_776
timestamp 1704896540
transform 1 0 72404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_782
timestamp 1704896540
transform 1 0 72956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_784
timestamp 1704896540
transform 1 0 73140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_796
timestamp 1704896540
transform 1 0 74244 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_800
timestamp 1704896540
transform 1 0 74612 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_702
timestamp 1704896540
transform 1 0 65596 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_714
timestamp 1704896540
transform 1 0 66700 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_726
timestamp 1704896540
transform 1 0 67804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_738
timestamp 1704896540
transform 1 0 68908 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_750
timestamp 1704896540
transform 1 0 70012 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_754
timestamp 1704896540
transform 1 0 70380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_756
timestamp 1704896540
transform 1 0 70564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_768
timestamp 1704896540
transform 1 0 71668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_780
timestamp 1704896540
transform 1 0 72772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_792
timestamp 1704896540
transform 1 0 73876 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_800
timestamp 1704896540
transform 1 0 74612 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_702
timestamp 1704896540
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_714
timestamp 1704896540
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_726
timestamp 1704896540
transform 1 0 67804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_728
timestamp 1704896540
transform 1 0 67988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_740
timestamp 1704896540
transform 1 0 69092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_752
timestamp 1704896540
transform 1 0 70196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_764
timestamp 1704896540
transform 1 0 71300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_776
timestamp 1704896540
transform 1 0 72404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_782
timestamp 1704896540
transform 1 0 72956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_784
timestamp 1704896540
transform 1 0 73140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_796
timestamp 1704896540
transform 1 0 74244 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_800
timestamp 1704896540
transform 1 0 74612 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_702
timestamp 1704896540
transform 1 0 65596 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_714
timestamp 1704896540
transform 1 0 66700 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_726
timestamp 1704896540
transform 1 0 67804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_738
timestamp 1704896540
transform 1 0 68908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_750
timestamp 1704896540
transform 1 0 70012 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_754
timestamp 1704896540
transform 1 0 70380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_756
timestamp 1704896540
transform 1 0 70564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_768
timestamp 1704896540
transform 1 0 71668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_780
timestamp 1704896540
transform 1 0 72772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_792
timestamp 1704896540
transform 1 0 73876 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_800
timestamp 1704896540
transform 1 0 74612 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_702
timestamp 1704896540
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_714
timestamp 1704896540
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_726
timestamp 1704896540
transform 1 0 67804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_728
timestamp 1704896540
transform 1 0 67988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_740
timestamp 1704896540
transform 1 0 69092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_752
timestamp 1704896540
transform 1 0 70196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_764
timestamp 1704896540
transform 1 0 71300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_776
timestamp 1704896540
transform 1 0 72404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_782
timestamp 1704896540
transform 1 0 72956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_784
timestamp 1704896540
transform 1 0 73140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_796
timestamp 1704896540
transform 1 0 74244 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_800
timestamp 1704896540
transform 1 0 74612 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_702
timestamp 1704896540
transform 1 0 65596 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_714
timestamp 1704896540
transform 1 0 66700 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_726
timestamp 1704896540
transform 1 0 67804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_738
timestamp 1704896540
transform 1 0 68908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_750
timestamp 1704896540
transform 1 0 70012 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_754
timestamp 1704896540
transform 1 0 70380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_756
timestamp 1704896540
transform 1 0 70564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_768
timestamp 1704896540
transform 1 0 71668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_780
timestamp 1704896540
transform 1 0 72772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_792
timestamp 1704896540
transform 1 0 73876 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_800
timestamp 1704896540
transform 1 0 74612 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_702
timestamp 1704896540
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_714
timestamp 1704896540
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_726
timestamp 1704896540
transform 1 0 67804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_728
timestamp 1704896540
transform 1 0 67988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_740
timestamp 1704896540
transform 1 0 69092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_752
timestamp 1704896540
transform 1 0 70196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_764
timestamp 1704896540
transform 1 0 71300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_776
timestamp 1704896540
transform 1 0 72404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_782
timestamp 1704896540
transform 1 0 72956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_784
timestamp 1704896540
transform 1 0 73140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_796
timestamp 1704896540
transform 1 0 74244 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_800
timestamp 1704896540
transform 1 0 74612 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_702
timestamp 1704896540
transform 1 0 65596 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_714
timestamp 1704896540
transform 1 0 66700 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_726
timestamp 1704896540
transform 1 0 67804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_738
timestamp 1704896540
transform 1 0 68908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_750
timestamp 1704896540
transform 1 0 70012 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_754
timestamp 1704896540
transform 1 0 70380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_756
timestamp 1704896540
transform 1 0 70564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_768
timestamp 1704896540
transform 1 0 71668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_780
timestamp 1704896540
transform 1 0 72772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_792
timestamp 1704896540
transform 1 0 73876 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_800
timestamp 1704896540
transform 1 0 74612 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_702
timestamp 1704896540
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_714
timestamp 1704896540
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_726
timestamp 1704896540
transform 1 0 67804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_728
timestamp 1704896540
transform 1 0 67988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_740
timestamp 1704896540
transform 1 0 69092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_752
timestamp 1704896540
transform 1 0 70196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_764
timestamp 1704896540
transform 1 0 71300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_776
timestamp 1704896540
transform 1 0 72404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_782
timestamp 1704896540
transform 1 0 72956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_784
timestamp 1704896540
transform 1 0 73140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_796
timestamp 1704896540
transform 1 0 74244 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_800
timestamp 1704896540
transform 1 0 74612 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_702
timestamp 1704896540
transform 1 0 65596 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_714
timestamp 1704896540
transform 1 0 66700 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_726
timestamp 1704896540
transform 1 0 67804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_738
timestamp 1704896540
transform 1 0 68908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_750
timestamp 1704896540
transform 1 0 70012 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_754
timestamp 1704896540
transform 1 0 70380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_756
timestamp 1704896540
transform 1 0 70564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_768
timestamp 1704896540
transform 1 0 71668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_780
timestamp 1704896540
transform 1 0 72772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_792
timestamp 1704896540
transform 1 0 73876 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_800
timestamp 1704896540
transform 1 0 74612 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_702
timestamp 1704896540
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_714
timestamp 1704896540
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_726
timestamp 1704896540
transform 1 0 67804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_728
timestamp 1704896540
transform 1 0 67988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_740
timestamp 1704896540
transform 1 0 69092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_752
timestamp 1704896540
transform 1 0 70196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_764
timestamp 1704896540
transform 1 0 71300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_776
timestamp 1704896540
transform 1 0 72404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_782
timestamp 1704896540
transform 1 0 72956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_784
timestamp 1704896540
transform 1 0 73140 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_796
timestamp 1704896540
transform 1 0 74244 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_800
timestamp 1704896540
transform 1 0 74612 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_702
timestamp 1704896540
transform 1 0 65596 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_714
timestamp 1704896540
transform 1 0 66700 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_726
timestamp 1704896540
transform 1 0 67804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_738
timestamp 1704896540
transform 1 0 68908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_750
timestamp 1704896540
transform 1 0 70012 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_754
timestamp 1704896540
transform 1 0 70380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_756
timestamp 1704896540
transform 1 0 70564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_768
timestamp 1704896540
transform 1 0 71668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_780
timestamp 1704896540
transform 1 0 72772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_792
timestamp 1704896540
transform 1 0 73876 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_800
timestamp 1704896540
transform 1 0 74612 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_702
timestamp 1704896540
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_714
timestamp 1704896540
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_726
timestamp 1704896540
transform 1 0 67804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_728
timestamp 1704896540
transform 1 0 67988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_740
timestamp 1704896540
transform 1 0 69092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_752
timestamp 1704896540
transform 1 0 70196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_764
timestamp 1704896540
transform 1 0 71300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_124_776
timestamp 1704896540
transform 1 0 72404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_782
timestamp 1704896540
transform 1 0 72956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_784
timestamp 1704896540
transform 1 0 73140 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124_796
timestamp 1704896540
transform 1 0 74244 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_800
timestamp 1704896540
transform 1 0 74612 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_702
timestamp 1704896540
transform 1 0 65596 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_714
timestamp 1704896540
transform 1 0 66700 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_726
timestamp 1704896540
transform 1 0 67804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_738
timestamp 1704896540
transform 1 0 68908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125_750
timestamp 1704896540
transform 1 0 70012 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_754
timestamp 1704896540
transform 1 0 70380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_756
timestamp 1704896540
transform 1 0 70564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_768
timestamp 1704896540
transform 1 0 71668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_780
timestamp 1704896540
transform 1 0 72772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_792
timestamp 1704896540
transform 1 0 73876 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_800
timestamp 1704896540
transform 1 0 74612 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_702
timestamp 1704896540
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_714
timestamp 1704896540
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_726
timestamp 1704896540
transform 1 0 67804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_728
timestamp 1704896540
transform 1 0 67988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_740
timestamp 1704896540
transform 1 0 69092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_752
timestamp 1704896540
transform 1 0 70196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_764
timestamp 1704896540
transform 1 0 71300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_126_776
timestamp 1704896540
transform 1 0 72404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_782
timestamp 1704896540
transform 1 0 72956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_784
timestamp 1704896540
transform 1 0 73140 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126_796
timestamp 1704896540
transform 1 0 74244 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_800
timestamp 1704896540
transform 1 0 74612 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_702
timestamp 1704896540
transform 1 0 65596 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_714
timestamp 1704896540
transform 1 0 66700 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_726
timestamp 1704896540
transform 1 0 67804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_738
timestamp 1704896540
transform 1 0 68908 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127_750
timestamp 1704896540
transform 1 0 70012 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_754
timestamp 1704896540
transform 1 0 70380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_756
timestamp 1704896540
transform 1 0 70564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_768
timestamp 1704896540
transform 1 0 71668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_780
timestamp 1704896540
transform 1 0 72772 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_792
timestamp 1704896540
transform 1 0 73876 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_800
timestamp 1704896540
transform 1 0 74612 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_702
timestamp 1704896540
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_714
timestamp 1704896540
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_726
timestamp 1704896540
transform 1 0 67804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_728
timestamp 1704896540
transform 1 0 67988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_740
timestamp 1704896540
transform 1 0 69092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_752
timestamp 1704896540
transform 1 0 70196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_764
timestamp 1704896540
transform 1 0 71300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_128_776
timestamp 1704896540
transform 1 0 72404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_782
timestamp 1704896540
transform 1 0 72956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_784
timestamp 1704896540
transform 1 0 73140 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128_796
timestamp 1704896540
transform 1 0 74244 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_800
timestamp 1704896540
transform 1 0 74612 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_702
timestamp 1704896540
transform 1 0 65596 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_714
timestamp 1704896540
transform 1 0 66700 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_726
timestamp 1704896540
transform 1 0 67804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_738
timestamp 1704896540
transform 1 0 68908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129_750
timestamp 1704896540
transform 1 0 70012 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_754
timestamp 1704896540
transform 1 0 70380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_756
timestamp 1704896540
transform 1 0 70564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_768
timestamp 1704896540
transform 1 0 71668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_780
timestamp 1704896540
transform 1 0 72772 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_792
timestamp 1704896540
transform 1 0 73876 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_800
timestamp 1704896540
transform 1 0 74612 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_702
timestamp 1704896540
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_714
timestamp 1704896540
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_726
timestamp 1704896540
transform 1 0 67804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_728
timestamp 1704896540
transform 1 0 67988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_740
timestamp 1704896540
transform 1 0 69092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_752
timestamp 1704896540
transform 1 0 70196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_764
timestamp 1704896540
transform 1 0 71300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_130_776
timestamp 1704896540
transform 1 0 72404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_782
timestamp 1704896540
transform 1 0 72956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_784
timestamp 1704896540
transform 1 0 73140 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130_796
timestamp 1704896540
transform 1 0 74244 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_800
timestamp 1704896540
transform 1 0 74612 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_702
timestamp 1704896540
transform 1 0 65596 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_714
timestamp 1704896540
transform 1 0 66700 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_726
timestamp 1704896540
transform 1 0 67804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_738
timestamp 1704896540
transform 1 0 68908 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131_750
timestamp 1704896540
transform 1 0 70012 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_754
timestamp 1704896540
transform 1 0 70380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_756
timestamp 1704896540
transform 1 0 70564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_768
timestamp 1704896540
transform 1 0 71668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_780
timestamp 1704896540
transform 1 0 72772 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_792
timestamp 1704896540
transform 1 0 73876 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_800
timestamp 1704896540
transform 1 0 74612 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_702
timestamp 1704896540
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_714
timestamp 1704896540
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_726
timestamp 1704896540
transform 1 0 67804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_728
timestamp 1704896540
transform 1 0 67988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_740
timestamp 1704896540
transform 1 0 69092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_752
timestamp 1704896540
transform 1 0 70196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_764
timestamp 1704896540
transform 1 0 71300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_132_776
timestamp 1704896540
transform 1 0 72404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_782
timestamp 1704896540
transform 1 0 72956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_784
timestamp 1704896540
transform 1 0 73140 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132_796
timestamp 1704896540
transform 1 0 74244 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_800
timestamp 1704896540
transform 1 0 74612 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_702
timestamp 1704896540
transform 1 0 65596 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_714
timestamp 1704896540
transform 1 0 66700 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_726
timestamp 1704896540
transform 1 0 67804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_738
timestamp 1704896540
transform 1 0 68908 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_750
timestamp 1704896540
transform 1 0 70012 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_754
timestamp 1704896540
transform 1 0 70380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_756
timestamp 1704896540
transform 1 0 70564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_768
timestamp 1704896540
transform 1 0 71668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_780
timestamp 1704896540
transform 1 0 72772 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_792
timestamp 1704896540
transform 1 0 73876 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_800
timestamp 1704896540
transform 1 0 74612 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_702
timestamp 1704896540
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_714
timestamp 1704896540
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_726
timestamp 1704896540
transform 1 0 67804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_728
timestamp 1704896540
transform 1 0 67988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_740
timestamp 1704896540
transform 1 0 69092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_752
timestamp 1704896540
transform 1 0 70196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_764
timestamp 1704896540
transform 1 0 71300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134_776
timestamp 1704896540
transform 1 0 72404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_782
timestamp 1704896540
transform 1 0 72956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_784
timestamp 1704896540
transform 1 0 73140 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134_796
timestamp 1704896540
transform 1 0 74244 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_800
timestamp 1704896540
transform 1 0 74612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_702
timestamp 1704896540
transform 1 0 65596 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_714
timestamp 1704896540
transform 1 0 66700 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_726
timestamp 1704896540
transform 1 0 67804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_738
timestamp 1704896540
transform 1 0 68908 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135_750
timestamp 1704896540
transform 1 0 70012 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_754
timestamp 1704896540
transform 1 0 70380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_756
timestamp 1704896540
transform 1 0 70564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_768
timestamp 1704896540
transform 1 0 71668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_780
timestamp 1704896540
transform 1 0 72772 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_792
timestamp 1704896540
transform 1 0 73876 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_800
timestamp 1704896540
transform 1 0 74612 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_702
timestamp 1704896540
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_714
timestamp 1704896540
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_726
timestamp 1704896540
transform 1 0 67804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_728
timestamp 1704896540
transform 1 0 67988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_740
timestamp 1704896540
transform 1 0 69092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_752
timestamp 1704896540
transform 1 0 70196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_764
timestamp 1704896540
transform 1 0 71300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_136_776
timestamp 1704896540
transform 1 0 72404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_782
timestamp 1704896540
transform 1 0 72956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_784
timestamp 1704896540
transform 1 0 73140 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136_796
timestamp 1704896540
transform 1 0 74244 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_800
timestamp 1704896540
transform 1 0 74612 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_702
timestamp 1704896540
transform 1 0 65596 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_714
timestamp 1704896540
transform 1 0 66700 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_726
timestamp 1704896540
transform 1 0 67804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_738
timestamp 1704896540
transform 1 0 68908 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137_750
timestamp 1704896540
transform 1 0 70012 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_754
timestamp 1704896540
transform 1 0 70380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_756
timestamp 1704896540
transform 1 0 70564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_768
timestamp 1704896540
transform 1 0 71668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_780
timestamp 1704896540
transform 1 0 72772 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_792
timestamp 1704896540
transform 1 0 73876 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_800
timestamp 1704896540
transform 1 0 74612 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_702
timestamp 1704896540
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_714
timestamp 1704896540
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_726
timestamp 1704896540
transform 1 0 67804 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_728
timestamp 1704896540
transform 1 0 67988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_740
timestamp 1704896540
transform 1 0 69092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_752
timestamp 1704896540
transform 1 0 70196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_764
timestamp 1704896540
transform 1 0 71300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_138_776
timestamp 1704896540
transform 1 0 72404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_782
timestamp 1704896540
transform 1 0 72956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_784
timestamp 1704896540
transform 1 0 73140 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_138_796
timestamp 1704896540
transform 1 0 74244 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_800
timestamp 1704896540
transform 1 0 74612 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_702
timestamp 1704896540
transform 1 0 65596 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_714
timestamp 1704896540
transform 1 0 66700 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_726
timestamp 1704896540
transform 1 0 67804 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_738
timestamp 1704896540
transform 1 0 68908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_139_750
timestamp 1704896540
transform 1 0 70012 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_754
timestamp 1704896540
transform 1 0 70380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_756
timestamp 1704896540
transform 1 0 70564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_768
timestamp 1704896540
transform 1 0 71668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_780
timestamp 1704896540
transform 1 0 72772 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_139_792
timestamp 1704896540
transform 1 0 73876 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_800
timestamp 1704896540
transform 1 0 74612 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_702
timestamp 1704896540
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_714
timestamp 1704896540
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_726
timestamp 1704896540
transform 1 0 67804 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_728
timestamp 1704896540
transform 1 0 67988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_740
timestamp 1704896540
transform 1 0 69092 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_752
timestamp 1704896540
transform 1 0 70196 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_764
timestamp 1704896540
transform 1 0 71300 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_140_776
timestamp 1704896540
transform 1 0 72404 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_782
timestamp 1704896540
transform 1 0 72956 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_784
timestamp 1704896540
transform 1 0 73140 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140_796
timestamp 1704896540
transform 1 0 74244 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_800
timestamp 1704896540
transform 1 0 74612 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_702
timestamp 1704896540
transform 1 0 65596 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_714
timestamp 1704896540
transform 1 0 66700 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_726
timestamp 1704896540
transform 1 0 67804 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_738
timestamp 1704896540
transform 1 0 68908 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141_750
timestamp 1704896540
transform 1 0 70012 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_754
timestamp 1704896540
transform 1 0 70380 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_756
timestamp 1704896540
transform 1 0 70564 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_768
timestamp 1704896540
transform 1 0 71668 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_780
timestamp 1704896540
transform 1 0 72772 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141_792
timestamp 1704896540
transform 1 0 73876 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_800
timestamp 1704896540
transform 1 0 74612 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_702
timestamp 1704896540
transform 1 0 65596 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_714
timestamp 1704896540
transform 1 0 66700 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_726
timestamp 1704896540
transform 1 0 67804 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_728
timestamp 1704896540
transform 1 0 67988 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_740
timestamp 1704896540
transform 1 0 69092 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_752
timestamp 1704896540
transform 1 0 70196 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_764
timestamp 1704896540
transform 1 0 71300 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_142_776
timestamp 1704896540
transform 1 0 72404 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_782
timestamp 1704896540
transform 1 0 72956 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_784
timestamp 1704896540
transform 1 0 73140 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142_796
timestamp 1704896540
transform 1 0 74244 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_800
timestamp 1704896540
transform 1 0 74612 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_702
timestamp 1704896540
transform 1 0 65596 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_714
timestamp 1704896540
transform 1 0 66700 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_726
timestamp 1704896540
transform 1 0 67804 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_738
timestamp 1704896540
transform 1 0 68908 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143_750
timestamp 1704896540
transform 1 0 70012 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_754
timestamp 1704896540
transform 1 0 70380 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_756
timestamp 1704896540
transform 1 0 70564 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_768
timestamp 1704896540
transform 1 0 71668 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_780
timestamp 1704896540
transform 1 0 72772 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_143_792
timestamp 1704896540
transform 1 0 73876 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_800
timestamp 1704896540
transform 1 0 74612 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_702
timestamp 1704896540
transform 1 0 65596 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_714
timestamp 1704896540
transform 1 0 66700 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_726
timestamp 1704896540
transform 1 0 67804 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_728
timestamp 1704896540
transform 1 0 67988 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_740
timestamp 1704896540
transform 1 0 69092 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_752
timestamp 1704896540
transform 1 0 70196 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_764
timestamp 1704896540
transform 1 0 71300 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144_776
timestamp 1704896540
transform 1 0 72404 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_782
timestamp 1704896540
transform 1 0 72956 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_784
timestamp 1704896540
transform 1 0 73140 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144_796
timestamp 1704896540
transform 1 0 74244 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_800
timestamp 1704896540
transform 1 0 74612 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_702
timestamp 1704896540
transform 1 0 65596 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_714
timestamp 1704896540
transform 1 0 66700 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_726
timestamp 1704896540
transform 1 0 67804 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_738
timestamp 1704896540
transform 1 0 68908 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145_750
timestamp 1704896540
transform 1 0 70012 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_754
timestamp 1704896540
transform 1 0 70380 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_756
timestamp 1704896540
transform 1 0 70564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_768
timestamp 1704896540
transform 1 0 71668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_780
timestamp 1704896540
transform 1 0 72772 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145_792
timestamp 1704896540
transform 1 0 73876 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_800
timestamp 1704896540
transform 1 0 74612 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_702
timestamp 1704896540
transform 1 0 65596 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_714
timestamp 1704896540
transform 1 0 66700 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_726
timestamp 1704896540
transform 1 0 67804 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_728
timestamp 1704896540
transform 1 0 67988 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_740
timestamp 1704896540
transform 1 0 69092 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_752
timestamp 1704896540
transform 1 0 70196 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_764
timestamp 1704896540
transform 1 0 71300 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146_776
timestamp 1704896540
transform 1 0 72404 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_782
timestamp 1704896540
transform 1 0 72956 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_784
timestamp 1704896540
transform 1 0 73140 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146_796
timestamp 1704896540
transform 1 0 74244 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_800
timestamp 1704896540
transform 1 0 74612 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_702
timestamp 1704896540
transform 1 0 65596 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_714
timestamp 1704896540
transform 1 0 66700 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_726
timestamp 1704896540
transform 1 0 67804 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_738
timestamp 1704896540
transform 1 0 68908 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147_750
timestamp 1704896540
transform 1 0 70012 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_754
timestamp 1704896540
transform 1 0 70380 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_756
timestamp 1704896540
transform 1 0 70564 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_768
timestamp 1704896540
transform 1 0 71668 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_780
timestamp 1704896540
transform 1 0 72772 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147_792
timestamp 1704896540
transform 1 0 73876 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_800
timestamp 1704896540
transform 1 0 74612 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_702
timestamp 1704896540
transform 1 0 65596 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_714
timestamp 1704896540
transform 1 0 66700 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_726
timestamp 1704896540
transform 1 0 67804 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_728
timestamp 1704896540
transform 1 0 67988 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_740
timestamp 1704896540
transform 1 0 69092 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_752
timestamp 1704896540
transform 1 0 70196 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_764
timestamp 1704896540
transform 1 0 71300 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_148_776
timestamp 1704896540
transform 1 0 72404 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_782
timestamp 1704896540
transform 1 0 72956 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_784
timestamp 1704896540
transform 1 0 73140 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148_796
timestamp 1704896540
transform 1 0 74244 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_800
timestamp 1704896540
transform 1 0 74612 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_702
timestamp 1704896540
transform 1 0 65596 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_714
timestamp 1704896540
transform 1 0 66700 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_726
timestamp 1704896540
transform 1 0 67804 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_738
timestamp 1704896540
transform 1 0 68908 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149_750
timestamp 1704896540
transform 1 0 70012 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_754
timestamp 1704896540
transform 1 0 70380 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_756
timestamp 1704896540
transform 1 0 70564 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_768
timestamp 1704896540
transform 1 0 71668 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_780
timestamp 1704896540
transform 1 0 72772 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_149_792
timestamp 1704896540
transform 1 0 73876 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_800
timestamp 1704896540
transform 1 0 74612 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_702
timestamp 1704896540
transform 1 0 65596 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_714
timestamp 1704896540
transform 1 0 66700 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_726
timestamp 1704896540
transform 1 0 67804 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_728
timestamp 1704896540
transform 1 0 67988 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_740
timestamp 1704896540
transform 1 0 69092 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_752
timestamp 1704896540
transform 1 0 70196 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_764
timestamp 1704896540
transform 1 0 71300 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_150_776
timestamp 1704896540
transform 1 0 72404 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_782
timestamp 1704896540
transform 1 0 72956 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_784
timestamp 1704896540
transform 1 0 73140 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150_796
timestamp 1704896540
transform 1 0 74244 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_800
timestamp 1704896540
transform 1 0 74612 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_702
timestamp 1704896540
transform 1 0 65596 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_714
timestamp 1704896540
transform 1 0 66700 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_726
timestamp 1704896540
transform 1 0 67804 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_738
timestamp 1704896540
transform 1 0 68908 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151_750
timestamp 1704896540
transform 1 0 70012 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_754
timestamp 1704896540
transform 1 0 70380 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_756
timestamp 1704896540
transform 1 0 70564 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_768
timestamp 1704896540
transform 1 0 71668 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_780
timestamp 1704896540
transform 1 0 72772 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151_792
timestamp 1704896540
transform 1 0 73876 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_800
timestamp 1704896540
transform 1 0 74612 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_702
timestamp 1704896540
transform 1 0 65596 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_714
timestamp 1704896540
transform 1 0 66700 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_726
timestamp 1704896540
transform 1 0 67804 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_728
timestamp 1704896540
transform 1 0 67988 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_740
timestamp 1704896540
transform 1 0 69092 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_752
timestamp 1704896540
transform 1 0 70196 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_764
timestamp 1704896540
transform 1 0 71300 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_152_776
timestamp 1704896540
transform 1 0 72404 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_782
timestamp 1704896540
transform 1 0 72956 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_784
timestamp 1704896540
transform 1 0 73140 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152_796
timestamp 1704896540
transform 1 0 74244 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_800
timestamp 1704896540
transform 1 0 74612 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_702
timestamp 1704896540
transform 1 0 65596 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_714
timestamp 1704896540
transform 1 0 66700 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_726
timestamp 1704896540
transform 1 0 67804 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_738
timestamp 1704896540
transform 1 0 68908 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153_750
timestamp 1704896540
transform 1 0 70012 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_754
timestamp 1704896540
transform 1 0 70380 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_756
timestamp 1704896540
transform 1 0 70564 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_768
timestamp 1704896540
transform 1 0 71668 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_780
timestamp 1704896540
transform 1 0 72772 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153_792
timestamp 1704896540
transform 1 0 73876 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_800
timestamp 1704896540
transform 1 0 74612 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_702
timestamp 1704896540
transform 1 0 65596 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_714
timestamp 1704896540
transform 1 0 66700 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_726
timestamp 1704896540
transform 1 0 67804 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_728
timestamp 1704896540
transform 1 0 67988 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_740
timestamp 1704896540
transform 1 0 69092 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_752
timestamp 1704896540
transform 1 0 70196 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_764
timestamp 1704896540
transform 1 0 71300 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154_776
timestamp 1704896540
transform 1 0 72404 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_782
timestamp 1704896540
transform 1 0 72956 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_784
timestamp 1704896540
transform 1 0 73140 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154_796
timestamp 1704896540
transform 1 0 74244 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_800
timestamp 1704896540
transform 1 0 74612 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_702
timestamp 1704896540
transform 1 0 65596 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_714
timestamp 1704896540
transform 1 0 66700 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_726
timestamp 1704896540
transform 1 0 67804 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_728
timestamp 1704896540
transform 1 0 67988 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_740
timestamp 1704896540
transform 1 0 69092 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_752
timestamp 1704896540
transform 1 0 70196 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_756
timestamp 1704896540
transform 1 0 70564 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_768
timestamp 1704896540
transform 1 0 71668 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_780
timestamp 1704896540
transform 1 0 72772 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_784
timestamp 1704896540
transform 1 0 73140 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_155_796
timestamp 1704896540
transform 1 0 74244 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_800
timestamp 1704896540
transform 1 0 74612 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 39836 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform 1 0 51244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 46092 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 55200 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 63756 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 66332 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 25208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform 1 0 44436 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform 1 0 21988 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform 1 0 43332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform 1 0 65964 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 66332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform 1 0 37444 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform 1 0 50416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 67988 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 66332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 45632 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform 1 0 54096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform 1 0 41952 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform 1 0 17480 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform 1 0 41216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 70012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform 1 0 36156 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform 1 0 49128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 44528 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform 1 0 53360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform 1 0 70932 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform 1 0 33948 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform 1 0 48944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 73968 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 68724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform 1 0 41032 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform 1 0 52624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform 1 0 32476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform 1 0 48208 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform 1 0 47472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform 1 0 28980 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform 1 0 47472 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform 1 0 53268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 66332 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform 1 0 51152 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 66332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform 1 0 49404 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 66332 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform -1 0 49680 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 66332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform 1 0 54372 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 66332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 57408 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 66332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform 1 0 59156 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 66332 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform 1 0 57776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform -1 0 66332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform -1 0 35972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 66332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 62560 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 66332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 27416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform 1 0 45356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform 1 0 62928 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 66332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform -1 0 66332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform 1 0 31188 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 66332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform 1 0 46368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform 1 0 26036 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform 1 0 45632 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform 1 0 44896 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 23184 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform 1 0 43792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform 1 0 19872 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform 1 0 17572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform 1 0 40388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold86 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 42964 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform 1 0 19136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold89
timestamp 1704896540
transform 1 0 42320 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold92
timestamp 1704896540
transform 1 0 65596 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold95
timestamp 1704896540
transform 1 0 65596 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform 1 0 24564 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform 1 0 43700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform -1 0 46184 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform -1 0 35880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform 1 0 29716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform 1 0 15732 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform -1 0 46920 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform -1 0 47104 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform -1 0 41952 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform -1 0 40572 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 37260 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform 1 0 34868 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform 1 0 33212 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1704896540
transform -1 0 33212 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1704896540
transform 1 0 29716 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1704896540
transform -1 0 54832 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1704896540
transform -1 0 52256 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1704896540
transform -1 0 30176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1704896540
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1704896540
transform 1 0 47380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1704896540
transform 1 0 54096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1704896540
transform -1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1704896540
transform -1 0 60076 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1704896540
transform 1 0 55476 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1704896540
transform -1 0 65136 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1704896540
transform 1 0 57316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1704896540
transform -1 0 28244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1704896540
transform 1 0 60444 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1704896540
transform -1 0 23920 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1704896540
transform 1 0 62284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1704896540
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1704896540
transform -1 0 68816 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1704896540
transform -1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1704896540
transform -1 0 19136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1704896540
transform 1 0 69552 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1704896540
transform 1 0 70656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1704896540
transform 1 0 72312 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1704896540
transform -1 0 36708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1704896540
transform 1 0 32292 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1704896540
transform -1 0 32476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1704896540
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1704896540
transform 1 0 27140 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1704896540
transform -1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1704896540
transform 1 0 23460 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1704896540
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1704896540
transform 1 0 16744 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform -1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1704896540
transform -1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 44528 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 47104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1704896540
transform -1 0 20240 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1704896540
transform -1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1704896540
transform -1 0 25300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1704896540
transform 1 0 26864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1704896540
transform -1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1704896540
transform -1 0 28980 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1704896540
transform 1 0 32016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1704896540
transform -1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1704896540
transform -1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform 1 0 16192 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input15
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1704896540
transform 1 0 38180 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1704896540
transform -1 0 39652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 41768 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1704896540
transform -1 0 42780 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1704896540
transform -1 0 44804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1704896540
transform 1 0 46920 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1704896540
transform -1 0 47380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1704896540
transform 1 0 50140 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1704896540
transform 1 0 51888 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1704896540
transform 1 0 54096 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1704896540
transform -1 0 19780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1704896540
transform 1 0 55200 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1704896540
transform -1 0 56304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1704896540
transform 1 0 58512 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1704896540
transform 1 0 59892 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1704896540
transform -1 0 61180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1704896540
transform -1 0 63572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1704896540
transform 1 0 65504 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1704896540
transform 1 0 66700 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1704896540
transform -1 0 67804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1704896540
transform -1 0 69460 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input37
timestamp 1704896540
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input38
timestamp 1704896540
transform 1 0 71668 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input39
timestamp 1704896540
transform -1 0 73140 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input40
timestamp 1704896540
transform -1 0 25852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1704896540
transform -1 0 27876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1704896540
transform -1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1704896540
transform -1 0 31740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1704896540
transform -1 0 33120 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1704896540
transform -1 0 34684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1704896540
transform -1 0 36432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input47
timestamp 1704896540
transform 1 0 19780 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input48
timestamp 1704896540
transform 1 0 21988 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input49
timestamp 1704896540
transform 1 0 24196 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input50
timestamp 1704896540
transform 1 0 26864 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1704896540
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18032 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1704896540
transform -1 0 5152 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1704896540
transform -1 0 18032 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1704896540
transform -1 0 21528 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1704896540
transform 1 0 37996 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1704896540
transform 1 0 39744 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1704896540
transform 1 0 42320 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1704896540
transform 1 0 42964 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1704896540
transform 1 0 44896 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1704896540
transform 1 0 47472 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1704896540
transform 1 0 47932 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1704896540
transform 1 0 50048 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1704896540
transform 1 0 52624 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1704896540
transform 1 0 52900 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1704896540
transform -1 0 22908 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1704896540
transform 1 0 55200 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1704896540
transform 1 0 56212 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1704896540
transform 1 0 57868 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1704896540
transform 1 0 60352 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1704896540
transform 1 0 61180 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1704896540
transform 1 0 62928 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1704896540
transform 1 0 64492 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1704896540
transform 1 0 66148 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1704896540
transform 1 0 68080 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1704896540
transform 1 0 69460 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1704896540
transform -1 0 24196 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1704896540
transform 1 0 71116 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1704896540
transform 1 0 73232 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1704896540
transform -1 0 26772 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1704896540
transform 1 0 27876 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1704896540
transform 1 0 29716 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1704896540
transform 1 0 30452 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1704896540
transform 1 0 33028 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1704896540
transform 1 0 34684 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1704896540
transform 1 0 35604 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_0
timestamp 1704896540
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_9
timestamp 1704896540
transform -1 0 74980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_1
timestamp 1704896540
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_10
timestamp 1704896540
transform -1 0 74980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_2
timestamp 1704896540
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_11
timestamp 1704896540
transform -1 0 74980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_3
timestamp 1704896540
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_12
timestamp 1704896540
transform -1 0 74980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_4
timestamp 1704896540
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_13
timestamp 1704896540
transform -1 0 74980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_5
timestamp 1704896540
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_14
timestamp 1704896540
transform -1 0 74980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_6
timestamp 1704896540
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_15
timestamp 1704896540
transform -1 0 74980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_7
timestamp 1704896540
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_16
timestamp 1704896540
transform -1 0 74980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_8
timestamp 1704896540
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_17
timestamp 1704896540
transform -1 0 74980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_311
timestamp 1704896540
transform 1 0 65320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_164
timestamp 1704896540
transform -1 0 74980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_165
timestamp 1704896540
transform 1 0 65320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_18
timestamp 1704896540
transform -1 0 74980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_166
timestamp 1704896540
transform 1 0 65320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_19
timestamp 1704896540
transform -1 0 74980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_167
timestamp 1704896540
transform 1 0 65320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_20
timestamp 1704896540
transform -1 0 74980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_168
timestamp 1704896540
transform 1 0 65320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_21
timestamp 1704896540
transform -1 0 74980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_169
timestamp 1704896540
transform 1 0 65320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_22
timestamp 1704896540
transform -1 0 74980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_170
timestamp 1704896540
transform 1 0 65320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_23
timestamp 1704896540
transform -1 0 74980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_171
timestamp 1704896540
transform 1 0 65320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_24
timestamp 1704896540
transform -1 0 74980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_172
timestamp 1704896540
transform 1 0 65320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_25
timestamp 1704896540
transform -1 0 74980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_173
timestamp 1704896540
transform 1 0 65320 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_26
timestamp 1704896540
transform -1 0 74980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_174
timestamp 1704896540
transform 1 0 65320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_27
timestamp 1704896540
transform -1 0 74980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_175
timestamp 1704896540
transform 1 0 65320 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_28
timestamp 1704896540
transform -1 0 74980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_176
timestamp 1704896540
transform 1 0 65320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_29
timestamp 1704896540
transform -1 0 74980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_177
timestamp 1704896540
transform 1 0 65320 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_30
timestamp 1704896540
transform -1 0 74980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_178
timestamp 1704896540
transform 1 0 65320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_31
timestamp 1704896540
transform -1 0 74980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_179
timestamp 1704896540
transform 1 0 65320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_32
timestamp 1704896540
transform -1 0 74980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_180
timestamp 1704896540
transform 1 0 65320 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_33
timestamp 1704896540
transform -1 0 74980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_181
timestamp 1704896540
transform 1 0 65320 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_34
timestamp 1704896540
transform -1 0 74980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_182
timestamp 1704896540
transform 1 0 65320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_35
timestamp 1704896540
transform -1 0 74980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_183
timestamp 1704896540
transform 1 0 65320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_36
timestamp 1704896540
transform -1 0 74980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_184
timestamp 1704896540
transform 1 0 65320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_37
timestamp 1704896540
transform -1 0 74980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_185
timestamp 1704896540
transform 1 0 65320 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_38
timestamp 1704896540
transform -1 0 74980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_186
timestamp 1704896540
transform 1 0 65320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_39
timestamp 1704896540
transform -1 0 74980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_187
timestamp 1704896540
transform 1 0 65320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_40
timestamp 1704896540
transform -1 0 74980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_188
timestamp 1704896540
transform 1 0 65320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_41
timestamp 1704896540
transform -1 0 74980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_189
timestamp 1704896540
transform 1 0 65320 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_42
timestamp 1704896540
transform -1 0 74980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_190
timestamp 1704896540
transform 1 0 65320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_43
timestamp 1704896540
transform -1 0 74980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_191
timestamp 1704896540
transform 1 0 65320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_44
timestamp 1704896540
transform -1 0 74980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_192
timestamp 1704896540
transform 1 0 65320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_45
timestamp 1704896540
transform -1 0 74980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_193
timestamp 1704896540
transform 1 0 65320 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_46
timestamp 1704896540
transform -1 0 74980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_194
timestamp 1704896540
transform 1 0 65320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_47
timestamp 1704896540
transform -1 0 74980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_195
timestamp 1704896540
transform 1 0 65320 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_48
timestamp 1704896540
transform -1 0 74980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_196
timestamp 1704896540
transform 1 0 65320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_49
timestamp 1704896540
transform -1 0 74980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_197
timestamp 1704896540
transform 1 0 65320 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_50
timestamp 1704896540
transform -1 0 74980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_198
timestamp 1704896540
transform 1 0 65320 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_51
timestamp 1704896540
transform -1 0 74980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_199
timestamp 1704896540
transform 1 0 65320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_52
timestamp 1704896540
transform -1 0 74980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_200
timestamp 1704896540
transform 1 0 65320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_53
timestamp 1704896540
transform -1 0 74980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_201
timestamp 1704896540
transform 1 0 65320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_54
timestamp 1704896540
transform -1 0 74980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_202
timestamp 1704896540
transform 1 0 65320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_55
timestamp 1704896540
transform -1 0 74980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_203
timestamp 1704896540
transform 1 0 65320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_56
timestamp 1704896540
transform -1 0 74980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_204
timestamp 1704896540
transform 1 0 65320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_57
timestamp 1704896540
transform -1 0 74980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_205
timestamp 1704896540
transform 1 0 65320 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_58
timestamp 1704896540
transform -1 0 74980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_206
timestamp 1704896540
transform 1 0 65320 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_59
timestamp 1704896540
transform -1 0 74980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_207
timestamp 1704896540
transform 1 0 65320 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_60
timestamp 1704896540
transform -1 0 74980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_208
timestamp 1704896540
transform 1 0 65320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_61
timestamp 1704896540
transform -1 0 74980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_209
timestamp 1704896540
transform 1 0 65320 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_62
timestamp 1704896540
transform -1 0 74980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_210
timestamp 1704896540
transform 1 0 65320 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_63
timestamp 1704896540
transform -1 0 74980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_211
timestamp 1704896540
transform 1 0 65320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_64
timestamp 1704896540
transform -1 0 74980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_212
timestamp 1704896540
transform 1 0 65320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_65
timestamp 1704896540
transform -1 0 74980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_213
timestamp 1704896540
transform 1 0 65320 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_66
timestamp 1704896540
transform -1 0 74980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_214
timestamp 1704896540
transform 1 0 65320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_67
timestamp 1704896540
transform -1 0 74980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_215
timestamp 1704896540
transform 1 0 65320 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_68
timestamp 1704896540
transform -1 0 74980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_216
timestamp 1704896540
transform 1 0 65320 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_69
timestamp 1704896540
transform -1 0 74980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_217
timestamp 1704896540
transform 1 0 65320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_70
timestamp 1704896540
transform -1 0 74980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_218
timestamp 1704896540
transform 1 0 65320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_71
timestamp 1704896540
transform -1 0 74980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_219
timestamp 1704896540
transform 1 0 65320 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_72
timestamp 1704896540
transform -1 0 74980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_220
timestamp 1704896540
transform 1 0 65320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_73
timestamp 1704896540
transform -1 0 74980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_221
timestamp 1704896540
transform 1 0 65320 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_74
timestamp 1704896540
transform -1 0 74980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_222
timestamp 1704896540
transform 1 0 65320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_75
timestamp 1704896540
transform -1 0 74980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_223
timestamp 1704896540
transform 1 0 65320 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_76
timestamp 1704896540
transform -1 0 74980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_224
timestamp 1704896540
transform 1 0 65320 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_77
timestamp 1704896540
transform -1 0 74980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_225
timestamp 1704896540
transform 1 0 65320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_78
timestamp 1704896540
transform -1 0 74980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_226
timestamp 1704896540
transform 1 0 65320 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_79
timestamp 1704896540
transform -1 0 74980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_227
timestamp 1704896540
transform 1 0 65320 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_80
timestamp 1704896540
transform -1 0 74980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_228
timestamp 1704896540
transform 1 0 65320 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_81
timestamp 1704896540
transform -1 0 74980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_229
timestamp 1704896540
transform 1 0 65320 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_82
timestamp 1704896540
transform -1 0 74980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_230
timestamp 1704896540
transform 1 0 65320 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_83
timestamp 1704896540
transform -1 0 74980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_231
timestamp 1704896540
transform 1 0 65320 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_84
timestamp 1704896540
transform -1 0 74980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_232
timestamp 1704896540
transform 1 0 65320 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_85
timestamp 1704896540
transform -1 0 74980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_233
timestamp 1704896540
transform 1 0 65320 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_86
timestamp 1704896540
transform -1 0 74980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_234
timestamp 1704896540
transform 1 0 65320 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_87
timestamp 1704896540
transform -1 0 74980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_235
timestamp 1704896540
transform 1 0 65320 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_88
timestamp 1704896540
transform -1 0 74980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_236
timestamp 1704896540
transform 1 0 65320 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_89
timestamp 1704896540
transform -1 0 74980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_237
timestamp 1704896540
transform 1 0 65320 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_90
timestamp 1704896540
transform -1 0 74980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_238
timestamp 1704896540
transform 1 0 65320 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_91
timestamp 1704896540
transform -1 0 74980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_239
timestamp 1704896540
transform 1 0 65320 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_92
timestamp 1704896540
transform -1 0 74980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_240
timestamp 1704896540
transform 1 0 65320 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_93
timestamp 1704896540
transform -1 0 74980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_241
timestamp 1704896540
transform 1 0 65320 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_94
timestamp 1704896540
transform -1 0 74980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_242
timestamp 1704896540
transform 1 0 65320 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_95
timestamp 1704896540
transform -1 0 74980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_243
timestamp 1704896540
transform 1 0 65320 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_96
timestamp 1704896540
transform -1 0 74980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_244
timestamp 1704896540
transform 1 0 65320 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_97
timestamp 1704896540
transform -1 0 74980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_245
timestamp 1704896540
transform 1 0 65320 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_98
timestamp 1704896540
transform -1 0 74980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_246
timestamp 1704896540
transform 1 0 65320 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_99
timestamp 1704896540
transform -1 0 74980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_247
timestamp 1704896540
transform 1 0 65320 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_100
timestamp 1704896540
transform -1 0 74980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_248
timestamp 1704896540
transform 1 0 65320 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_101
timestamp 1704896540
transform -1 0 74980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_249
timestamp 1704896540
transform 1 0 65320 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_102
timestamp 1704896540
transform -1 0 74980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_250
timestamp 1704896540
transform 1 0 65320 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_103
timestamp 1704896540
transform -1 0 74980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_251
timestamp 1704896540
transform 1 0 65320 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_104
timestamp 1704896540
transform -1 0 74980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_252
timestamp 1704896540
transform 1 0 65320 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_105
timestamp 1704896540
transform -1 0 74980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_253
timestamp 1704896540
transform 1 0 65320 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_106
timestamp 1704896540
transform -1 0 74980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_254
timestamp 1704896540
transform 1 0 65320 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_107
timestamp 1704896540
transform -1 0 74980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_255
timestamp 1704896540
transform 1 0 65320 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_108
timestamp 1704896540
transform -1 0 74980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_256
timestamp 1704896540
transform 1 0 65320 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_109
timestamp 1704896540
transform -1 0 74980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_257
timestamp 1704896540
transform 1 0 65320 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_110
timestamp 1704896540
transform -1 0 74980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_258
timestamp 1704896540
transform 1 0 65320 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_111
timestamp 1704896540
transform -1 0 74980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_259
timestamp 1704896540
transform 1 0 65320 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_112
timestamp 1704896540
transform -1 0 74980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_260
timestamp 1704896540
transform 1 0 65320 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_113
timestamp 1704896540
transform -1 0 74980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_261
timestamp 1704896540
transform 1 0 65320 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_114
timestamp 1704896540
transform -1 0 74980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_262
timestamp 1704896540
transform 1 0 65320 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_115
timestamp 1704896540
transform -1 0 74980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_263
timestamp 1704896540
transform 1 0 65320 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_116
timestamp 1704896540
transform -1 0 74980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_264
timestamp 1704896540
transform 1 0 65320 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_117
timestamp 1704896540
transform -1 0 74980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_265
timestamp 1704896540
transform 1 0 65320 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_118
timestamp 1704896540
transform -1 0 74980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_266
timestamp 1704896540
transform 1 0 65320 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_119
timestamp 1704896540
transform -1 0 74980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_267
timestamp 1704896540
transform 1 0 65320 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_120
timestamp 1704896540
transform -1 0 74980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_268
timestamp 1704896540
transform 1 0 65320 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_121
timestamp 1704896540
transform -1 0 74980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_269
timestamp 1704896540
transform 1 0 65320 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_122
timestamp 1704896540
transform -1 0 74980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_270
timestamp 1704896540
transform 1 0 65320 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_123
timestamp 1704896540
transform -1 0 74980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_271
timestamp 1704896540
transform 1 0 65320 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_124
timestamp 1704896540
transform -1 0 74980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Left_272
timestamp 1704896540
transform 1 0 65320 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Right_125
timestamp 1704896540
transform -1 0 74980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Left_273
timestamp 1704896540
transform 1 0 65320 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Right_126
timestamp 1704896540
transform -1 0 74980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Left_274
timestamp 1704896540
transform 1 0 65320 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Right_127
timestamp 1704896540
transform -1 0 74980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Left_275
timestamp 1704896540
transform 1 0 65320 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Right_128
timestamp 1704896540
transform -1 0 74980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_276
timestamp 1704896540
transform 1 0 65320 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_129
timestamp 1704896540
transform -1 0 74980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_277
timestamp 1704896540
transform 1 0 65320 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_130
timestamp 1704896540
transform -1 0 74980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_278
timestamp 1704896540
transform 1 0 65320 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_131
timestamp 1704896540
transform -1 0 74980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_279
timestamp 1704896540
transform 1 0 65320 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_132
timestamp 1704896540
transform -1 0 74980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_280
timestamp 1704896540
transform 1 0 65320 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_133
timestamp 1704896540
transform -1 0 74980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_281
timestamp 1704896540
transform 1 0 65320 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_134
timestamp 1704896540
transform -1 0 74980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_282
timestamp 1704896540
transform 1 0 65320 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_135
timestamp 1704896540
transform -1 0 74980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_283
timestamp 1704896540
transform 1 0 65320 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_136
timestamp 1704896540
transform -1 0 74980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_284
timestamp 1704896540
transform 1 0 65320 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_137
timestamp 1704896540
transform -1 0 74980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_285
timestamp 1704896540
transform 1 0 65320 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_138
timestamp 1704896540
transform -1 0 74980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_286
timestamp 1704896540
transform 1 0 65320 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_139
timestamp 1704896540
transform -1 0 74980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_287
timestamp 1704896540
transform 1 0 65320 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_140
timestamp 1704896540
transform -1 0 74980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_288
timestamp 1704896540
transform 1 0 65320 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_141
timestamp 1704896540
transform -1 0 74980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_289
timestamp 1704896540
transform 1 0 65320 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_142
timestamp 1704896540
transform -1 0 74980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_290
timestamp 1704896540
transform 1 0 65320 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_143
timestamp 1704896540
transform -1 0 74980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_291
timestamp 1704896540
transform 1 0 65320 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_144
timestamp 1704896540
transform -1 0 74980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_292
timestamp 1704896540
transform 1 0 65320 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_145
timestamp 1704896540
transform -1 0 74980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_293
timestamp 1704896540
transform 1 0 65320 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_146
timestamp 1704896540
transform -1 0 74980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_294
timestamp 1704896540
transform 1 0 65320 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_147
timestamp 1704896540
transform -1 0 74980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_295
timestamp 1704896540
transform 1 0 65320 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_148
timestamp 1704896540
transform -1 0 74980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_296
timestamp 1704896540
transform 1 0 65320 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_149
timestamp 1704896540
transform -1 0 74980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_297
timestamp 1704896540
transform 1 0 65320 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_150
timestamp 1704896540
transform -1 0 74980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_298
timestamp 1704896540
transform 1 0 65320 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_151
timestamp 1704896540
transform -1 0 74980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_299
timestamp 1704896540
transform 1 0 65320 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_152
timestamp 1704896540
transform -1 0 74980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_300
timestamp 1704896540
transform 1 0 65320 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_153
timestamp 1704896540
transform -1 0 74980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_301
timestamp 1704896540
transform 1 0 65320 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_154
timestamp 1704896540
transform -1 0 74980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_302
timestamp 1704896540
transform 1 0 65320 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_155
timestamp 1704896540
transform -1 0 74980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_303
timestamp 1704896540
transform 1 0 65320 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_156
timestamp 1704896540
transform -1 0 74980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_304
timestamp 1704896540
transform 1 0 65320 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_157
timestamp 1704896540
transform -1 0 74980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_305
timestamp 1704896540
transform 1 0 65320 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_158
timestamp 1704896540
transform -1 0 74980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_306
timestamp 1704896540
transform 1 0 65320 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_159
timestamp 1704896540
transform -1 0 74980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_307
timestamp 1704896540
transform 1 0 65320 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_160
timestamp 1704896540
transform -1 0 74980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_308
timestamp 1704896540
transform 1 0 65320 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_161
timestamp 1704896540
transform -1 0 74980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_309
timestamp 1704896540
transform 1 0 65320 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_162
timestamp 1704896540
transform -1 0 74980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_310
timestamp 1704896540
transform 1 0 65320 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_163
timestamp 1704896540
transform -1 0 74980 0 -1 85952
box -38 -48 314 592
use EFSRAM_1024x32_wrapper  SRAM_0
timestamp 0
transform 0 -1 63283 1 0 8000
box 0 -40 77574 61263
use sky130_fd_sc_hd__conb_1  SRAM_0_87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 65872 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_88
timestamp 1704896540
transform -1 0 65872 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_89
timestamp 1704896540
transform -1 0 65872 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_90
timestamp 1704896540
transform -1 0 65872 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_91
timestamp 1704896540
transform -1 0 65872 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_92
timestamp 1704896540
transform -1 0 66148 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_93
timestamp 1704896540
transform -1 0 65872 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_94
timestamp 1704896540
transform 1 0 65596 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_95
timestamp 1704896540
transform 1 0 65872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_312 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_313
timestamp 1704896540
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_314
timestamp 1704896540
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_315
timestamp 1704896540
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_316
timestamp 1704896540
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_317
timestamp 1704896540
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_318
timestamp 1704896540
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_319
timestamp 1704896540
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_320
timestamp 1704896540
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_321
timestamp 1704896540
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_322
timestamp 1704896540
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_323
timestamp 1704896540
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_324
timestamp 1704896540
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_325
timestamp 1704896540
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_326
timestamp 1704896540
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_327
timestamp 1704896540
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_328
timestamp 1704896540
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_329
timestamp 1704896540
transform 1 0 47380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_330
timestamp 1704896540
transform 1 0 49956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_331
timestamp 1704896540
transform 1 0 52532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_332
timestamp 1704896540
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_333
timestamp 1704896540
transform 1 0 57684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_334
timestamp 1704896540
transform 1 0 60260 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_335
timestamp 1704896540
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_336
timestamp 1704896540
transform 1 0 65412 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_337
timestamp 1704896540
transform 1 0 67988 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_338
timestamp 1704896540
transform 1 0 70564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_339
timestamp 1704896540
transform 1 0 73140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_340
timestamp 1704896540
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_341
timestamp 1704896540
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_342
timestamp 1704896540
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_343
timestamp 1704896540
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_344
timestamp 1704896540
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_345
timestamp 1704896540
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_346
timestamp 1704896540
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_347
timestamp 1704896540
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_348
timestamp 1704896540
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_349
timestamp 1704896540
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_350
timestamp 1704896540
transform 1 0 57684 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_351
timestamp 1704896540
transform 1 0 62836 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_352
timestamp 1704896540
transform 1 0 67988 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_353
timestamp 1704896540
transform 1 0 73140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_354
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_355
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_356
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_357
timestamp 1704896540
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_358
timestamp 1704896540
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_359
timestamp 1704896540
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_360
timestamp 1704896540
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_361
timestamp 1704896540
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_362
timestamp 1704896540
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_363
timestamp 1704896540
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_364
timestamp 1704896540
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_365
timestamp 1704896540
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_366
timestamp 1704896540
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_367
timestamp 1704896540
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_368
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_369
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_370
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_371
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_372
timestamp 1704896540
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_373
timestamp 1704896540
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_374
timestamp 1704896540
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_375
timestamp 1704896540
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_376
timestamp 1704896540
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_377
timestamp 1704896540
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_378
timestamp 1704896540
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_379
timestamp 1704896540
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_380
timestamp 1704896540
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_381
timestamp 1704896540
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_382
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_383
timestamp 1704896540
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_384
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_385
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_386
timestamp 1704896540
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_387
timestamp 1704896540
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_388
timestamp 1704896540
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_389
timestamp 1704896540
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_390
timestamp 1704896540
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_391
timestamp 1704896540
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_392
timestamp 1704896540
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_393
timestamp 1704896540
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_394
timestamp 1704896540
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_395
timestamp 1704896540
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_396
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_397
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_398
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_399
timestamp 1704896540
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_400
timestamp 1704896540
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_401
timestamp 1704896540
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_402
timestamp 1704896540
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_403
timestamp 1704896540
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_404
timestamp 1704896540
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_405
timestamp 1704896540
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_406
timestamp 1704896540
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_407
timestamp 1704896540
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_408
timestamp 1704896540
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_409
timestamp 1704896540
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_410
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_411
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_412
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_413
timestamp 1704896540
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_414
timestamp 1704896540
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_415
timestamp 1704896540
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_416
timestamp 1704896540
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_417
timestamp 1704896540
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_418
timestamp 1704896540
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_419
timestamp 1704896540
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_420
timestamp 1704896540
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_421
timestamp 1704896540
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_422
timestamp 1704896540
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_423
timestamp 1704896540
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_424
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_425
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_426
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_427
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_428
timestamp 1704896540
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_429
timestamp 1704896540
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_430
timestamp 1704896540
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_431
timestamp 1704896540
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_432
timestamp 1704896540
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_433
timestamp 1704896540
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_434
timestamp 1704896540
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_435
timestamp 1704896540
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_436
timestamp 1704896540
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_437
timestamp 1704896540
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_438
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_439
timestamp 1704896540
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_440
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_441
timestamp 1704896540
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_442
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_443
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_444
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_445
timestamp 1704896540
transform 1 0 21620 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_446
timestamp 1704896540
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_447
timestamp 1704896540
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_448
timestamp 1704896540
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_449
timestamp 1704896540
transform 1 0 31924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_450
timestamp 1704896540
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_451
timestamp 1704896540
transform 1 0 37076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_452
timestamp 1704896540
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_453
timestamp 1704896540
transform 1 0 42228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_454
timestamp 1704896540
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_455
timestamp 1704896540
transform 1 0 47380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_456
timestamp 1704896540
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_457
timestamp 1704896540
transform 1 0 52532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_458
timestamp 1704896540
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_459
timestamp 1704896540
transform 1 0 57684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_460
timestamp 1704896540
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_461
timestamp 1704896540
transform 1 0 62836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_462
timestamp 1704896540
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_463
timestamp 1704896540
transform 1 0 67988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_464
timestamp 1704896540
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_465
timestamp 1704896540
transform 1 0 73140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_687
timestamp 1704896540
transform 1 0 70472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_466
timestamp 1704896540
transform 1 0 67896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_467
timestamp 1704896540
transform 1 0 73048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_468
timestamp 1704896540
transform 1 0 70472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_469
timestamp 1704896540
transform 1 0 67896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_470
timestamp 1704896540
transform 1 0 73048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_471
timestamp 1704896540
transform 1 0 70472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_472
timestamp 1704896540
transform 1 0 67896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_473
timestamp 1704896540
transform 1 0 73048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_474
timestamp 1704896540
transform 1 0 70472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_475
timestamp 1704896540
transform 1 0 67896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_476
timestamp 1704896540
transform 1 0 73048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_477
timestamp 1704896540
transform 1 0 70472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_478
timestamp 1704896540
transform 1 0 67896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_479
timestamp 1704896540
transform 1 0 73048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_480
timestamp 1704896540
transform 1 0 70472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_481
timestamp 1704896540
transform 1 0 67896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_482
timestamp 1704896540
transform 1 0 73048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_483
timestamp 1704896540
transform 1 0 70472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_484
timestamp 1704896540
transform 1 0 67896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_485
timestamp 1704896540
transform 1 0 73048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_486
timestamp 1704896540
transform 1 0 70472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_487
timestamp 1704896540
transform 1 0 67896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_488
timestamp 1704896540
transform 1 0 73048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_489
timestamp 1704896540
transform 1 0 70472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_490
timestamp 1704896540
transform 1 0 67896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_491
timestamp 1704896540
transform 1 0 73048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_492
timestamp 1704896540
transform 1 0 70472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_493
timestamp 1704896540
transform 1 0 67896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_494
timestamp 1704896540
transform 1 0 73048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_495
timestamp 1704896540
transform 1 0 70472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_496
timestamp 1704896540
transform 1 0 67896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_497
timestamp 1704896540
transform 1 0 73048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_498
timestamp 1704896540
transform 1 0 70472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_499
timestamp 1704896540
transform 1 0 67896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_500
timestamp 1704896540
transform 1 0 73048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_501
timestamp 1704896540
transform 1 0 70472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_502
timestamp 1704896540
transform 1 0 67896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_503
timestamp 1704896540
transform 1 0 73048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_504
timestamp 1704896540
transform 1 0 70472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_505
timestamp 1704896540
transform 1 0 67896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_506
timestamp 1704896540
transform 1 0 73048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_507
timestamp 1704896540
transform 1 0 70472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_508
timestamp 1704896540
transform 1 0 67896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_509
timestamp 1704896540
transform 1 0 73048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_510
timestamp 1704896540
transform 1 0 70472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_511
timestamp 1704896540
transform 1 0 67896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_512
timestamp 1704896540
transform 1 0 73048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_513
timestamp 1704896540
transform 1 0 70472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_514
timestamp 1704896540
transform 1 0 67896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_515
timestamp 1704896540
transform 1 0 73048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_516
timestamp 1704896540
transform 1 0 70472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_517
timestamp 1704896540
transform 1 0 67896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_518
timestamp 1704896540
transform 1 0 73048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_519
timestamp 1704896540
transform 1 0 70472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_520
timestamp 1704896540
transform 1 0 67896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_521
timestamp 1704896540
transform 1 0 73048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_522
timestamp 1704896540
transform 1 0 70472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_523
timestamp 1704896540
transform 1 0 67896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_524
timestamp 1704896540
transform 1 0 73048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_525
timestamp 1704896540
transform 1 0 70472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_526
timestamp 1704896540
transform 1 0 67896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_527
timestamp 1704896540
transform 1 0 73048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_528
timestamp 1704896540
transform 1 0 70472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_529
timestamp 1704896540
transform 1 0 67896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_530
timestamp 1704896540
transform 1 0 73048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_531
timestamp 1704896540
transform 1 0 70472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_532
timestamp 1704896540
transform 1 0 67896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_533
timestamp 1704896540
transform 1 0 73048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_534
timestamp 1704896540
transform 1 0 70472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_535
timestamp 1704896540
transform 1 0 67896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_536
timestamp 1704896540
transform 1 0 73048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_537
timestamp 1704896540
transform 1 0 70472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_538
timestamp 1704896540
transform 1 0 67896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_539
timestamp 1704896540
transform 1 0 73048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_540
timestamp 1704896540
transform 1 0 70472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_541
timestamp 1704896540
transform 1 0 67896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_542
timestamp 1704896540
transform 1 0 73048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_543
timestamp 1704896540
transform 1 0 70472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_544
timestamp 1704896540
transform 1 0 67896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_545
timestamp 1704896540
transform 1 0 73048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_546
timestamp 1704896540
transform 1 0 70472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_547
timestamp 1704896540
transform 1 0 67896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_548
timestamp 1704896540
transform 1 0 73048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_549
timestamp 1704896540
transform 1 0 70472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_550
timestamp 1704896540
transform 1 0 67896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_551
timestamp 1704896540
transform 1 0 73048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_552
timestamp 1704896540
transform 1 0 70472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_553
timestamp 1704896540
transform 1 0 67896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_554
timestamp 1704896540
transform 1 0 73048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_555
timestamp 1704896540
transform 1 0 70472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_556
timestamp 1704896540
transform 1 0 67896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_557
timestamp 1704896540
transform 1 0 73048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_558
timestamp 1704896540
transform 1 0 70472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_559
timestamp 1704896540
transform 1 0 67896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_560
timestamp 1704896540
transform 1 0 73048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_561
timestamp 1704896540
transform 1 0 70472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_562
timestamp 1704896540
transform 1 0 67896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_563
timestamp 1704896540
transform 1 0 73048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_564
timestamp 1704896540
transform 1 0 70472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_565
timestamp 1704896540
transform 1 0 67896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_566
timestamp 1704896540
transform 1 0 73048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_567
timestamp 1704896540
transform 1 0 70472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_568
timestamp 1704896540
transform 1 0 67896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_569
timestamp 1704896540
transform 1 0 73048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_570
timestamp 1704896540
transform 1 0 70472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_571
timestamp 1704896540
transform 1 0 67896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_572
timestamp 1704896540
transform 1 0 73048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_573
timestamp 1704896540
transform 1 0 70472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_574
timestamp 1704896540
transform 1 0 67896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_575
timestamp 1704896540
transform 1 0 73048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_576
timestamp 1704896540
transform 1 0 70472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_577
timestamp 1704896540
transform 1 0 67896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_578
timestamp 1704896540
transform 1 0 73048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_579
timestamp 1704896540
transform 1 0 70472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_580
timestamp 1704896540
transform 1 0 67896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_581
timestamp 1704896540
transform 1 0 73048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_582
timestamp 1704896540
transform 1 0 70472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_583
timestamp 1704896540
transform 1 0 67896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_584
timestamp 1704896540
transform 1 0 73048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_585
timestamp 1704896540
transform 1 0 70472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_586
timestamp 1704896540
transform 1 0 67896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_587
timestamp 1704896540
transform 1 0 73048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_588
timestamp 1704896540
transform 1 0 70472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_589
timestamp 1704896540
transform 1 0 67896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_590
timestamp 1704896540
transform 1 0 73048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_591
timestamp 1704896540
transform 1 0 70472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_592
timestamp 1704896540
transform 1 0 67896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_593
timestamp 1704896540
transform 1 0 73048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_594
timestamp 1704896540
transform 1 0 70472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_595
timestamp 1704896540
transform 1 0 67896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_596
timestamp 1704896540
transform 1 0 73048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_597
timestamp 1704896540
transform 1 0 70472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_598
timestamp 1704896540
transform 1 0 67896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_599
timestamp 1704896540
transform 1 0 73048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_600
timestamp 1704896540
transform 1 0 70472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_601
timestamp 1704896540
transform 1 0 67896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_602
timestamp 1704896540
transform 1 0 73048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_603
timestamp 1704896540
transform 1 0 70472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_604
timestamp 1704896540
transform 1 0 67896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_605
timestamp 1704896540
transform 1 0 73048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_606
timestamp 1704896540
transform 1 0 70472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_607
timestamp 1704896540
transform 1 0 67896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_608
timestamp 1704896540
transform 1 0 73048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_609
timestamp 1704896540
transform 1 0 70472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_610
timestamp 1704896540
transform 1 0 67896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_611
timestamp 1704896540
transform 1 0 73048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_612
timestamp 1704896540
transform 1 0 70472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_613
timestamp 1704896540
transform 1 0 67896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_614
timestamp 1704896540
transform 1 0 73048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_615
timestamp 1704896540
transform 1 0 70472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_616
timestamp 1704896540
transform 1 0 67896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_617
timestamp 1704896540
transform 1 0 73048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_618
timestamp 1704896540
transform 1 0 70472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_619
timestamp 1704896540
transform 1 0 67896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_620
timestamp 1704896540
transform 1 0 73048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_621
timestamp 1704896540
transform 1 0 70472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_622
timestamp 1704896540
transform 1 0 67896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_623
timestamp 1704896540
transform 1 0 73048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_624
timestamp 1704896540
transform 1 0 70472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_625
timestamp 1704896540
transform 1 0 67896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_626
timestamp 1704896540
transform 1 0 73048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_627
timestamp 1704896540
transform 1 0 70472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_628
timestamp 1704896540
transform 1 0 67896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_629
timestamp 1704896540
transform 1 0 73048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_630
timestamp 1704896540
transform 1 0 70472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_631
timestamp 1704896540
transform 1 0 67896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_632
timestamp 1704896540
transform 1 0 73048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_633
timestamp 1704896540
transform 1 0 70472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_634
timestamp 1704896540
transform 1 0 67896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_635
timestamp 1704896540
transform 1 0 73048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_636
timestamp 1704896540
transform 1 0 70472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_637
timestamp 1704896540
transform 1 0 67896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_638
timestamp 1704896540
transform 1 0 73048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_639
timestamp 1704896540
transform 1 0 70472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_640
timestamp 1704896540
transform 1 0 67896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_641
timestamp 1704896540
transform 1 0 73048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_642
timestamp 1704896540
transform 1 0 70472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_643
timestamp 1704896540
transform 1 0 67896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_644
timestamp 1704896540
transform 1 0 73048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_645
timestamp 1704896540
transform 1 0 70472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_646
timestamp 1704896540
transform 1 0 67896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_647
timestamp 1704896540
transform 1 0 73048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_648
timestamp 1704896540
transform 1 0 70472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_649
timestamp 1704896540
transform 1 0 67896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_650
timestamp 1704896540
transform 1 0 73048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_651
timestamp 1704896540
transform 1 0 70472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_652
timestamp 1704896540
transform 1 0 67896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_653
timestamp 1704896540
transform 1 0 73048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_654
timestamp 1704896540
transform 1 0 70472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_655
timestamp 1704896540
transform 1 0 67896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_656
timestamp 1704896540
transform 1 0 73048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_657
timestamp 1704896540
transform 1 0 70472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_658
timestamp 1704896540
transform 1 0 67896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_659
timestamp 1704896540
transform 1 0 73048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_660
timestamp 1704896540
transform 1 0 70472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_661
timestamp 1704896540
transform 1 0 67896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_662
timestamp 1704896540
transform 1 0 73048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_663
timestamp 1704896540
transform 1 0 70472 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_664
timestamp 1704896540
transform 1 0 67896 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_665
timestamp 1704896540
transform 1 0 73048 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_666
timestamp 1704896540
transform 1 0 70472 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_667
timestamp 1704896540
transform 1 0 67896 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_668
timestamp 1704896540
transform 1 0 73048 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_669
timestamp 1704896540
transform 1 0 70472 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_670
timestamp 1704896540
transform 1 0 67896 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_671
timestamp 1704896540
transform 1 0 73048 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_672
timestamp 1704896540
transform 1 0 70472 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_673
timestamp 1704896540
transform 1 0 67896 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_674
timestamp 1704896540
transform 1 0 73048 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_675
timestamp 1704896540
transform 1 0 70472 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_676
timestamp 1704896540
transform 1 0 67896 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_677
timestamp 1704896540
transform 1 0 73048 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_678
timestamp 1704896540
transform 1 0 70472 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_679
timestamp 1704896540
transform 1 0 67896 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_680
timestamp 1704896540
transform 1 0 73048 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_681
timestamp 1704896540
transform 1 0 70472 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_682
timestamp 1704896540
transform 1 0 67896 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_683
timestamp 1704896540
transform 1 0 73048 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_684
timestamp 1704896540
transform 1 0 67896 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_685
timestamp 1704896540
transform 1 0 70472 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_686
timestamp 1704896540
transform 1 0 73048 0 -1 85952
box -38 -48 130 592
<< labels >>
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 sram_selected
port 0 nsew signal tristate
flabel metal2 s 1836 1040 2188 5944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 11836 1040 12188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 21836 1040 22188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 31836 1040 32188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 41836 1040 42188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 51836 1040 52188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 61836 1040 62188 5972 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 71836 1040 72188 86000 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 1912 75028 2264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 11912 75028 12264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 21912 75028 22264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 31912 75028 32264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 41912 75028 42264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 51912 75028 52264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 61912 75028 62264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 71912 75028 72264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 964 81912 75028 82264 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 1702 86940 2322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 7702 86940 8322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 13702 86940 14322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 19702 86940 20322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 25702 86940 26322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 31702 86940 32322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 37702 86940 38322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 43702 86940 44322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 49702 86940 50322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 55702 86940 56322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 61702 86940 62322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 67702 86940 68322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 87000 0 FreeSans 3840 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 60 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal4 s 73702 86940 74322 87000 0 FreeSans 480 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 4188 1040 4540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 14188 1040 14540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 24188 1040 24540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 34188 1040 34540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 44188 1040 44540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 54188 1040 54540 5944 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 64188 1040 64540 5972 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 74188 1040 74540 86000 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 4264 75028 4616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 14264 75028 14616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 24264 75028 24616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 34264 75028 34616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 44264 75028 44616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 54264 75028 54616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 64264 75028 64616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 74264 75028 74616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 964 84264 75028 84616 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 0 5322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 0 5322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 4702 86940 5322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 0 11322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 0 11322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 10702 86940 11322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 0 17322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 0 17322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 16702 86940 17322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 0 23322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 0 23322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 22702 86940 23322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 0 29322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 0 29322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 28702 86940 29322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 0 35322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 0 35322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 34702 86940 35322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 0 41322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 0 41322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 40702 86940 41322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 0 47322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 0 47322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 46702 86940 47322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 0 53322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 0 53322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 52702 86940 53322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 0 59322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 0 59322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 58702 86940 59322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 0 65322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 0 65322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 64702 86940 65322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 0 71322 87000 0 FreeSans 3840 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 0 71322 60 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal4 s 70702 86940 71322 87000 0 FreeSans 480 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wb_clk_i
port 3 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wb_rst_i
port 4 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 5 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 6 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 7 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 8 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 9 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 10 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 11 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 12 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 13 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 14 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 15 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 16 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 17 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 18 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 19 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 20 nsew signal input
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 21 nsew signal input
flabel metal2 s 60002 0 60058 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 22 nsew signal input
flabel metal2 s 61658 0 61714 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 23 nsew signal input
flabel metal2 s 63314 0 63370 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 24 nsew signal input
flabel metal2 s 64970 0 65026 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 25 nsew signal input
flabel metal2 s 66626 0 66682 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 26 nsew signal input
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 27 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 28 nsew signal input
flabel metal2 s 69938 0 69994 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 29 nsew signal input
flabel metal2 s 71594 0 71650 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 30 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 31 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 32 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 33 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 34 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 35 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 36 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 37 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 38 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 39 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 40 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 41 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 42 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 43 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 44 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 45 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 46 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 47 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 48 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 49 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 50 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 51 nsew signal input
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 52 nsew signal input
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 53 nsew signal input
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 54 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 55 nsew signal input
flabel metal2 s 62210 0 62266 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 56 nsew signal input
flabel metal2 s 63866 0 63922 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 57 nsew signal input
flabel metal2 s 65522 0 65578 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 58 nsew signal input
flabel metal2 s 67178 0 67234 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 59 nsew signal input
flabel metal2 s 68834 0 68890 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 60 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 61 nsew signal input
flabel metal2 s 70490 0 70546 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 62 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 63 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 64 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 65 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 66 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 67 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 68 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 69 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 70 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 71 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 72 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 73 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 74 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 75 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 76 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 77 nsew signal tristate
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 78 nsew signal tristate
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 79 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 80 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 81 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 82 nsew signal tristate
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 83 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 84 nsew signal tristate
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 85 nsew signal tristate
flabel metal2 s 59450 0 59506 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 86 nsew signal tristate
flabel metal2 s 61106 0 61162 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 87 nsew signal tristate
flabel metal2 s 62762 0 62818 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 88 nsew signal tristate
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 89 nsew signal tristate
flabel metal2 s 66074 0 66130 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 90 nsew signal tristate
flabel metal2 s 67730 0 67786 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 91 nsew signal tristate
flabel metal2 s 69386 0 69442 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 92 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 93 nsew signal tristate
flabel metal2 s 71042 0 71098 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 94 nsew signal tristate
flabel metal2 s 72698 0 72754 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 95 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 96 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 97 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 98 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 99 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 100 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 101 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 102 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 103 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 104 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 105 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 106 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 107 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_we_i
port 108 nsew signal input
rlabel via2 62434 82208 62434 82208 0 vccd1
rlabel via2 62636 84560 62636 84560 0 vssd1
rlabel metal1 19826 1870 19826 1870 0 _000_
rlabel metal1 19327 2006 19327 2006 0 _001_
rlabel metal2 31694 4522 31694 4522 0 _002_
rlabel metal2 32246 4624 32246 4624 0 _003_
rlabel metal2 32338 4930 32338 4930 0 _004_
rlabel metal2 33350 4454 33350 4454 0 _005_
rlabel metal2 34914 4658 34914 4658 0 _006_
rlabel metal2 36846 4182 36846 4182 0 _007_
rlabel metal2 45954 3740 45954 3740 0 _008_
rlabel metal1 47334 3026 47334 3026 0 _009_
rlabel metal2 49082 3740 49082 3740 0 _010_
rlabel metal1 65642 5678 65642 5678 0 _011_
rlabel metal2 52946 4012 52946 4012 0 _012_
rlabel metal2 54694 4012 54694 4012 0 _013_
rlabel metal2 56258 4420 56258 4420 0 _014_
rlabel metal2 57822 4386 57822 4386 0 _015_
rlabel metal2 59478 4284 59478 4284 0 _016_
rlabel metal2 61226 4284 61226 4284 0 _017_
rlabel metal2 63250 4284 63250 4284 0 _018_
rlabel metal2 64814 4284 64814 4284 0 _019_
rlabel metal2 66470 4284 66470 4284 0 _020_
rlabel metal2 68126 4284 68126 4284 0 _021_
rlabel metal2 69874 4012 69874 4012 0 _022_
rlabel metal2 71438 4012 71438 4012 0 _023_
rlabel metal1 73094 3026 73094 3026 0 _024_
rlabel metal1 17526 2482 17526 2482 0 _025_
rlabel metal1 28014 3706 28014 3706 0 _026_
rlabel metal2 24886 4182 24886 4182 0 _027_
rlabel metal1 72588 5202 72588 5202 0 _028_
rlabel metal1 28198 2550 28198 2550 0 _029_
rlabel metal1 26404 3026 26404 3026 0 _030_
rlabel metal1 26726 3060 26726 3060 0 _031_
rlabel metal1 28428 3502 28428 3502 0 _032_
rlabel metal2 28566 4012 28566 4012 0 _033_
rlabel metal1 28336 2414 28336 2414 0 _034_
rlabel metal2 29486 2043 29486 2043 0 _035_
rlabel metal2 30038 3910 30038 3910 0 _036_
rlabel metal1 29716 3026 29716 3026 0 _037_
rlabel metal2 34730 4318 34730 4318 0 _038_
rlabel metal2 31234 4386 31234 4386 0 _039_
rlabel metal3 67091 33252 67091 33252 0 clknet_0_wb_clk_i
rlabel metal1 35834 5542 35834 5542 0 clknet_1_0__leaf_wb_clk_i
rlabel metal1 63250 53280 63250 53280 0 clknet_1_1__leaf_wb_clk_i
rlabel metal2 20746 1972 20746 1972 0 net1
rlabel metal2 36202 2346 36202 2346 0 net10
rlabel metal2 65182 1530 65182 1530 0 net100
rlabel metal1 63250 72262 63250 72262 0 net101
rlabel metal1 25852 3162 25852 3162 0 net102
rlabel metal1 63250 36405 63250 36405 0 net103
rlabel metal1 22816 1530 22816 1530 0 net104
rlabel metal1 63250 38699 63250 38699 0 net105
rlabel metal1 66700 1938 66700 1938 0 net106
rlabel metal1 63250 74590 63250 74590 0 net107
rlabel metal1 38226 1938 38226 1938 0 net108
rlabel metal1 63250 21159 63250 21159 0 net109
rlabel via3 66539 23460 66539 23460 0 net11
rlabel metal2 67298 2244 67298 2244 0 net110
rlabel metal1 63250 76618 63250 76618 0 net111
rlabel metal1 44850 2414 44850 2414 0 net112
rlabel metal1 63250 12563 63250 12563 0 net113
rlabel metal2 20286 3910 20286 3910 0 net114
rlabel metal1 63395 40838 63395 40838 0 net115
rlabel metal1 18216 2074 18216 2074 0 net116
rlabel metal1 63395 43018 63395 43018 0 net117
rlabel metal2 69414 2108 69414 2108 0 net118
rlabel metal1 63250 78796 63250 78796 0 net119
rlabel metal1 66424 23086 66424 23086 0 net12
rlabel metal1 36800 2074 36800 2074 0 net120
rlabel metal1 63250 23337 63250 23337 0 net121
rlabel metal1 43378 1326 43378 1326 0 net122
rlabel metal1 63250 14625 63250 14625 0 net123
rlabel metal1 71668 1938 71668 1938 0 net124
rlabel metal1 63250 81008 63250 81008 0 net125
rlabel metal1 34592 3026 34592 3026 0 net126
rlabel metal1 63250 25413 63250 25413 0 net127
rlabel metal1 73140 1326 73140 1326 0 net128
rlabel metal1 63250 83186 63250 83186 0 net129
rlabel metal1 39054 2380 39054 2380 0 net13
rlabel metal1 41768 1938 41768 1938 0 net130
rlabel metal1 63250 16735 63250 16735 0 net131
rlabel metal1 33074 3026 33074 3026 0 net132
rlabel metal1 63250 27693 63250 27693 0 net133
rlabel metal1 31648 2618 31648 2618 0 net134
rlabel metal1 63250 29769 63250 29769 0 net135
rlabel metal1 29624 1938 29624 1938 0 net136
rlabel metal1 63250 31947 63250 31947 0 net137
rlabel metal1 54096 3026 54096 3026 0 net138
rlabel metal1 63250 57016 63250 57016 0 net139
rlabel metal2 18354 2142 18354 2142 0 net14
rlabel metal1 51934 1938 51934 1938 0 net140
rlabel metal1 63250 54872 63250 54872 0 net141
rlabel metal1 50186 1938 50186 1938 0 net142
rlabel metal1 63250 52660 63250 52660 0 net143
rlabel metal1 48944 1326 48944 1326 0 net144
rlabel metal1 63250 50516 63250 50516 0 net145
rlabel metal2 55062 2210 55062 2210 0 net146
rlabel metal1 63250 59194 63250 59194 0 net147
rlabel metal2 56718 1836 56718 1836 0 net148
rlabel metal1 63250 61372 63250 61372 0 net149
rlabel metal2 41262 4114 41262 4114 0 net15
rlabel metal1 59938 1938 59938 1938 0 net150
rlabel metal1 63250 65728 63250 65728 0 net151
rlabel metal1 58558 1938 58558 1938 0 net152
rlabel metal1 63250 63584 63250 63584 0 net153
rlabel metal1 35236 2414 35236 2414 0 net154
rlabel metal1 63250 44445 63250 44445 0 net155
rlabel metal1 61456 1530 61456 1530 0 net156
rlabel metal1 63250 67906 63250 67906 0 net157
rlabel metal1 27922 3162 27922 3162 0 net158
rlabel metal1 63250 34125 63250 34125 0 net159
rlabel metal2 38594 1598 38594 1598 0 net16
rlabel metal2 63618 2210 63618 2210 0 net160
rlabel metal1 63250 70084 63250 70084 0 net161
rlabel metal1 34178 2618 34178 2618 0 net162
rlabel metal1 63618 44526 63618 44526 0 net163
rlabel metal1 32108 2074 32108 2074 0 net164
rlabel metal1 63250 45003 63250 45003 0 net165
rlabel metal1 28934 1904 28934 1904 0 net166
rlabel metal1 63802 45254 63802 45254 0 net167
rlabel metal1 29210 2618 29210 2618 0 net168
rlabel metal1 63710 45730 63710 45730 0 net169
rlabel metal2 39330 2312 39330 2312 0 net17
rlabel metal1 26864 2074 26864 2074 0 net170
rlabel metal1 63848 45934 63848 45934 0 net171
rlabel metal2 25254 3060 25254 3060 0 net172
rlabel metal1 63756 43826 63756 43826 0 net173
rlabel metal1 19734 1292 19734 1292 0 net174
rlabel metal1 63572 47022 63572 47022 0 net175
rlabel metal2 20562 3332 20562 3332 0 net176
rlabel metal1 64124 47362 64124 47362 0 net177
rlabel metal1 18216 2618 18216 2618 0 net178
rlabel via3 64469 47668 64469 47668 0 net179
rlabel metal2 52670 4658 52670 4658 0 net18
rlabel metal1 22310 1938 22310 1938 0 net180
rlabel metal1 63250 22271 63250 22271 0 net181
rlabel metal1 21574 2618 21574 2618 0 net182
rlabel metal2 19826 2074 19826 2074 0 net183
rlabel metal1 63250 37517 63250 37517 0 net184
rlabel metal1 19090 2618 19090 2618 0 net185
rlabel metal1 24702 1938 24702 1938 0 net186
rlabel metal1 63158 60274 63158 60274 0 net187
rlabel metal1 24104 2618 24104 2618 0 net188
rlabel metal1 26818 1938 26818 1938 0 net189
rlabel metal2 53406 3706 53406 3706 0 net19
rlabel metal1 63250 81904 63250 81904 0 net190
rlabel metal1 25668 1530 25668 1530 0 net191
rlabel metal1 44666 1326 44666 1326 0 net192
rlabel metal1 44758 1904 44758 1904 0 net193
rlabel metal1 32614 2856 32614 2856 0 net194
rlabel metal2 33994 4250 33994 4250 0 net195
rlabel metal1 18078 1258 18078 1258 0 net196
rlabel metal2 46230 2142 46230 2142 0 net197
rlabel metal1 46000 1530 46000 1530 0 net198
rlabel metal1 44482 1360 44482 1360 0 net199
rlabel metal2 17894 3536 17894 3536 0 net2
rlabel metal1 54326 3978 54326 3978 0 net20
rlabel metal1 41216 1530 41216 1530 0 net200
rlabel metal1 39836 1870 39836 1870 0 net201
rlabel metal1 37766 1530 37766 1530 0 net202
rlabel metal2 36202 1564 36202 1564 0 net203
rlabel metal1 33948 1870 33948 1870 0 net204
rlabel metal2 32522 2244 32522 2244 0 net205
rlabel metal1 30728 1530 30728 1530 0 net206
rlabel metal1 54004 1326 54004 1326 0 net207
rlabel metal1 51428 1530 51428 1530 0 net208
rlabel metal2 29118 2108 29118 2108 0 net209
rlabel metal2 55338 4114 55338 4114 0 net21
rlabel metal2 49542 2108 49542 2108 0 net210
rlabel metal1 49496 1326 49496 1326 0 net211
rlabel metal1 54648 1938 54648 1938 0 net212
rlabel metal2 25346 2788 25346 2788 0 net213
rlabel metal2 59386 1598 59386 1598 0 net214
rlabel metal2 57270 1530 57270 1530 0 net215
rlabel metal1 64170 1530 64170 1530 0 net216
rlabel metal2 57914 2108 57914 2108 0 net217
rlabel metal2 27554 2788 27554 2788 0 net218
rlabel metal2 62422 1530 62422 1530 0 net219
rlabel metal1 66792 23766 66792 23766 0 net22
rlabel metal1 22310 1326 22310 1326 0 net220
rlabel metal2 62974 2108 62974 2108 0 net221
rlabel metal2 66102 2108 66102 2108 0 net222
rlabel metal1 68034 1870 68034 1870 0 net223
rlabel metal1 20424 2618 20424 2618 0 net224
rlabel metal1 18032 1938 18032 1938 0 net225
rlabel metal1 70104 1530 70104 1530 0 net226
rlabel metal2 71070 2108 71070 2108 0 net227
rlabel metal1 73416 1870 73416 1870 0 net228
rlabel metal1 35972 2414 35972 2414 0 net229
rlabel metal3 66631 23324 66631 23324 0 net23
rlabel metal1 33304 1190 33304 1190 0 net230
rlabel metal2 31326 2108 31326 2108 0 net231
rlabel metal2 30958 2720 30958 2720 0 net232
rlabel metal1 28244 1530 28244 1530 0 net233
rlabel metal1 26174 1972 26174 1972 0 net234
rlabel metal1 24380 2074 24380 2074 0 net235
rlabel metal2 23138 3196 23138 3196 0 net236
rlabel metal2 19918 2788 19918 2788 0 net237
rlabel metal1 17526 2074 17526 2074 0 net238
rlabel metal1 54050 1802 54050 1802 0 net24
rlabel metal1 66378 29614 66378 29614 0 net25
rlabel metal1 27738 4080 27738 4080 0 net26
rlabel metal1 63066 2312 63066 2312 0 net27
rlabel metal1 58420 2618 58420 2618 0 net28
rlabel metal1 60030 2074 60030 2074 0 net29
rlabel metal1 45402 1190 45402 1190 0 net3
rlabel metal2 65458 2159 65458 2159 0 net30
rlabel metal1 63296 2482 63296 2482 0 net31
rlabel metal1 65366 2618 65366 2618 0 net32
rlabel metal1 65826 1224 65826 1224 0 net33
rlabel metal1 66976 2006 66976 2006 0 net34
rlabel metal1 66884 39406 66884 39406 0 net35
rlabel metal1 69184 2006 69184 2006 0 net36
rlabel metal1 31878 2312 31878 2312 0 net37
rlabel metal1 71070 2006 71070 2006 0 net38
rlabel metal1 71438 1258 71438 1258 0 net39
rlabel metal1 47058 1530 47058 1530 0 net4
rlabel metal2 28842 3519 28842 3519 0 net40
rlabel metal2 33074 4590 33074 4590 0 net41
rlabel metal1 29532 3162 29532 3162 0 net42
rlabel metal2 33442 3434 33442 3434 0 net43
rlabel metal2 32614 4386 32614 4386 0 net44
rlabel metal1 34086 2822 34086 2822 0 net45
rlabel metal1 35972 3094 35972 3094 0 net46
rlabel metal1 21551 1394 21551 1394 0 net47
rlabel metal2 41722 4964 41722 4964 0 net48
rlabel metal1 60030 2516 60030 2516 0 net49
rlabel metal2 40618 4930 40618 4930 0 net5
rlabel metal1 64860 2040 64860 2040 0 net50
rlabel metal1 21252 2958 21252 2958 0 net51
rlabel metal1 20378 4148 20378 4148 0 net52
rlabel metal2 5106 1156 5106 1156 0 net53
rlabel metal2 17802 1802 17802 1802 0 net54
rlabel metal1 21482 1972 21482 1972 0 net55
rlabel metal1 35558 3502 35558 3502 0 net56
rlabel metal2 39790 2448 39790 2448 0 net57
rlabel metal2 36938 3196 36938 3196 0 net58
rlabel metal1 35650 3060 35650 3060 0 net59
rlabel metal2 19458 1054 19458 1054 0 net6
rlabel metal1 35098 2856 35098 2856 0 net60
rlabel metal2 37030 3264 37030 3264 0 net61
rlabel metal1 47794 1938 47794 1938 0 net62
rlabel metal1 48898 2890 48898 2890 0 net63
rlabel metal2 52670 2074 52670 2074 0 net64
rlabel metal2 53130 2380 53130 2380 0 net65
rlabel metal1 22862 2448 22862 2448 0 net66
rlabel metal1 55062 2822 55062 2822 0 net67
rlabel metal2 56442 2380 56442 2380 0 net68
rlabel metal2 58006 2074 58006 2074 0 net69
rlabel metal2 24978 4862 24978 4862 0 net7
rlabel metal1 60030 2822 60030 2822 0 net70
rlabel metal2 61410 2380 61410 2380 0 net71
rlabel metal2 63066 2074 63066 2074 0 net72
rlabel metal2 64630 2380 64630 2380 0 net73
rlabel metal2 66286 2074 66286 2074 0 net74
rlabel metal2 68310 2074 68310 2074 0 net75
rlabel metal2 69690 2380 69690 2380 0 net76
rlabel metal1 24150 1258 24150 1258 0 net77
rlabel metal2 71254 2074 71254 2074 0 net78
rlabel metal2 73278 2074 73278 2074 0 net79
rlabel metal2 27094 4590 27094 4590 0 net8
rlabel metal1 26726 1258 26726 1258 0 net80
rlabel metal1 28244 2822 28244 2822 0 net81
rlabel metal1 29762 1972 29762 1972 0 net82
rlabel metal1 30498 1292 30498 1292 0 net83
rlabel metal2 33258 2210 33258 2210 0 net84
rlabel metal1 32522 2924 32522 2924 0 net85
rlabel metal2 35650 1156 35650 1156 0 net86
rlabel metal1 63618 49631 63618 49631 0 net87
rlabel metal1 63250 43713 63250 43713 0 net88
rlabel metal1 63250 42543 63250 42543 0 net89
rlabel metal2 28658 4726 28658 4726 0 net9
rlabel metal1 63250 50114 63250 50114 0 net90
rlabel metal1 63441 52094 63441 52094 0 net91
rlabel metal1 63250 52289 63250 52289 0 net92
rlabel metal1 63441 48715 63441 48715 0 net93
rlabel metal1 67022 47022 67022 47022 0 net94
rlabel metal1 66562 46954 66562 46954 0 net95
rlabel metal2 39146 2210 39146 2210 0 net96
rlabel metal1 63250 18879 63250 18879 0 net97
rlabel metal1 46920 1938 46920 1938 0 net98
rlabel metal1 56028 5678 56028 5678 0 net99
rlabel metal1 63250 43283 63250 43283 0 ram_controller.DO\[0\]
rlabel metal1 63441 21470 63441 21470 0 ram_controller.DO\[10\]
rlabel metal1 63250 19209 63250 19209 0 ram_controller.DO\[11\]
rlabel metal1 63441 17110 63441 17110 0 ram_controller.DO\[12\]
rlabel metal1 63250 14853 63250 14853 0 ram_controller.DO\[13\]
rlabel metal1 64085 12750 64085 12750 0 ram_controller.DO\[14\]
rlabel metal2 27554 5950 27554 5950 0 ram_controller.DO\[15\]
rlabel metal1 63250 50288 63250 50288 0 ram_controller.DO\[16\]
rlabel metal1 63158 52466 63158 52466 0 ram_controller.DO\[17\]
rlabel metal1 63250 54576 63250 54576 0 ram_controller.DO\[18\]
rlabel metal1 63441 56844 63441 56844 0 ram_controller.DO\[19\]
rlabel metal1 63250 41023 63250 41023 0 ram_controller.DO\[1\]
rlabel metal1 63250 59048 63250 59048 0 ram_controller.DO\[20\]
rlabel metal1 63250 61042 63250 61042 0 ram_controller.DO\[21\]
rlabel metal1 63250 63288 63250 63288 0 ram_controller.DO\[22\]
rlabel metal1 63250 65582 63250 65582 0 ram_controller.DO\[23\]
rlabel metal1 63395 67744 63395 67744 0 ram_controller.DO\[24\]
rlabel metal3 63365 17884 63365 17884 0 ram_controller.DO\[25\]
rlabel metal1 63250 71932 63250 71932 0 ram_controller.DO\[26\]
rlabel metal1 63250 74178 63250 74178 0 ram_controller.DO\[27\]
rlabel metal1 63250 76472 63250 76472 0 ram_controller.DO\[28\]
rlabel metal1 63250 78636 63250 78636 0 ram_controller.DO\[29\]
rlabel metal1 63250 38845 63250 38845 0 ram_controller.DO\[2\]
rlabel metal1 63250 80814 63250 80814 0 ram_controller.DO\[30\]
rlabel metal1 63250 82992 63250 82992 0 ram_controller.DO\[31\]
rlabel metal1 63250 36633 63250 36633 0 ram_controller.DO\[3\]
rlabel metal1 63441 34550 63441 34550 0 ram_controller.DO\[4\]
rlabel metal1 63250 32277 63250 32277 0 ram_controller.DO\[5\]
rlabel metal1 63250 30099 63250 30099 0 ram_controller.DO\[6\]
rlabel metal1 63250 27921 63250 27921 0 ram_controller.DO\[7\]
rlabel metal1 63250 25743 63250 25743 0 ram_controller.DO\[8\]
rlabel metal1 63250 23565 63250 23565 0 ram_controller.DO\[9\]
rlabel metal1 63250 48969 63250 48969 0 ram_controller.EN
rlabel metal1 63250 48105 63250 48105 0 ram_controller.R_WB
rlabel metal2 20654 3298 20654 3298 0 ram_controller.wbs_ack_o
rlabel metal2 3174 1010 3174 1010 0 sram_selected
rlabel metal2 14766 2047 14766 2047 0 wb_clk_i
rlabel metal2 15318 1044 15318 1044 0 wb_rst_i
rlabel metal2 15870 823 15870 823 0 wbs_ack_o
rlabel metal2 18078 1316 18078 1316 0 wbs_adr_i[0]
rlabel metal2 43470 1588 43470 1588 0 wbs_adr_i[14]
rlabel metal2 45126 1010 45126 1010 0 wbs_adr_i[15]
rlabel metal2 20286 1588 20286 1588 0 wbs_adr_i[1]
rlabel metal1 22540 3502 22540 3502 0 wbs_adr_i[2]
rlabel metal2 24702 1316 24702 1316 0 wbs_adr_i[3]
rlabel metal2 26910 1588 26910 1588 0 wbs_adr_i[4]
rlabel metal2 28566 1010 28566 1010 0 wbs_adr_i[5]
rlabel metal1 30268 2958 30268 2958 0 wbs_adr_i[6]
rlabel metal2 31878 823 31878 823 0 wbs_adr_i[7]
rlabel metal2 33534 840 33534 840 0 wbs_adr_i[8]
rlabel metal2 36570 1938 36570 1938 0 wbs_adr_i[9]
rlabel metal2 16422 1350 16422 1350 0 wbs_cyc_i
rlabel metal2 18630 1163 18630 1163 0 wbs_dat_i[0]
rlabel metal2 37398 1044 37398 1044 0 wbs_dat_i[10]
rlabel metal2 39054 1350 39054 1350 0 wbs_dat_i[11]
rlabel metal2 40710 1044 40710 1044 0 wbs_dat_i[12]
rlabel metal2 42366 1588 42366 1588 0 wbs_dat_i[13]
rlabel metal2 44022 1010 44022 1010 0 wbs_dat_i[14]
rlabel metal2 45678 1350 45678 1350 0 wbs_dat_i[15]
rlabel metal2 47334 1588 47334 1588 0 wbs_dat_i[16]
rlabel metal2 48990 1588 48990 1588 0 wbs_dat_i[17]
rlabel metal2 50646 1044 50646 1044 0 wbs_dat_i[18]
rlabel metal2 52302 976 52302 976 0 wbs_dat_i[19]
rlabel metal2 20838 1622 20838 1622 0 wbs_dat_i[1]
rlabel metal2 53958 1588 53958 1588 0 wbs_dat_i[20]
rlabel metal2 55614 1316 55614 1316 0 wbs_dat_i[21]
rlabel metal2 57270 959 57270 959 0 wbs_dat_i[22]
rlabel metal2 58926 1010 58926 1010 0 wbs_dat_i[23]
rlabel metal2 60582 1316 60582 1316 0 wbs_dat_i[24]
rlabel metal2 62238 1027 62238 1027 0 wbs_dat_i[25]
rlabel metal2 63894 1044 63894 1044 0 wbs_dat_i[26]
rlabel metal2 65550 1588 65550 1588 0 wbs_dat_i[27]
rlabel metal2 67206 1350 67206 1350 0 wbs_dat_i[28]
rlabel metal2 68862 1044 68862 1044 0 wbs_dat_i[29]
rlabel metal1 23414 2958 23414 2958 0 wbs_dat_i[2]
rlabel metal2 70518 1588 70518 1588 0 wbs_dat_i[30]
rlabel metal2 72174 823 72174 823 0 wbs_dat_i[31]
rlabel metal2 25254 1588 25254 1588 0 wbs_dat_i[3]
rlabel metal2 27462 1588 27462 1588 0 wbs_dat_i[4]
rlabel metal2 29118 1027 29118 1027 0 wbs_dat_i[5]
rlabel metal2 30774 823 30774 823 0 wbs_dat_i[6]
rlabel metal2 32430 1316 32430 1316 0 wbs_dat_i[7]
rlabel metal2 34086 1350 34086 1350 0 wbs_dat_i[8]
rlabel metal2 35742 976 35742 976 0 wbs_dat_i[9]
rlabel metal2 19182 1095 19182 1095 0 wbs_dat_o[0]
rlabel metal2 37950 1078 37950 1078 0 wbs_dat_o[10]
rlabel metal2 39606 1010 39606 1010 0 wbs_dat_o[11]
rlabel metal2 41262 1078 41262 1078 0 wbs_dat_o[12]
rlabel metal2 42918 891 42918 891 0 wbs_dat_o[13]
rlabel metal2 44574 823 44574 823 0 wbs_dat_o[14]
rlabel metal2 46230 1078 46230 1078 0 wbs_dat_o[15]
rlabel metal2 47886 1316 47886 1316 0 wbs_dat_o[16]
rlabel metal2 49542 1078 49542 1078 0 wbs_dat_o[17]
rlabel metal2 51198 1010 51198 1010 0 wbs_dat_o[18]
rlabel metal2 52854 1316 52854 1316 0 wbs_dat_o[19]
rlabel metal2 21390 1588 21390 1588 0 wbs_dat_o[1]
rlabel metal2 54510 823 54510 823 0 wbs_dat_o[20]
rlabel metal2 56166 1316 56166 1316 0 wbs_dat_o[21]
rlabel metal2 57822 1010 57822 1010 0 wbs_dat_o[22]
rlabel metal2 59478 1078 59478 1078 0 wbs_dat_o[23]
rlabel metal2 61134 1316 61134 1316 0 wbs_dat_o[24]
rlabel metal2 62790 1078 62790 1078 0 wbs_dat_o[25]
rlabel metal2 64446 823 64446 823 0 wbs_dat_o[26]
rlabel metal2 66102 1010 66102 1010 0 wbs_dat_o[27]
rlabel metal2 67758 1078 67758 1078 0 wbs_dat_o[28]
rlabel metal2 69414 1282 69414 1282 0 wbs_dat_o[29]
rlabel metal2 23598 1010 23598 1010 0 wbs_dat_o[2]
rlabel metal2 71070 1078 71070 1078 0 wbs_dat_o[30]
rlabel metal2 72726 976 72726 976 0 wbs_dat_o[31]
rlabel metal2 25806 1010 25806 1010 0 wbs_dat_o[3]
rlabel metal2 28014 1078 28014 1078 0 wbs_dat_o[4]
rlabel metal2 29670 823 29670 823 0 wbs_dat_o[5]
rlabel metal2 31326 1010 31326 1010 0 wbs_dat_o[6]
rlabel metal2 32982 1010 32982 1010 0 wbs_dat_o[7]
rlabel metal2 34638 1316 34638 1316 0 wbs_dat_o[8]
rlabel metal2 36294 1010 36294 1010 0 wbs_dat_o[9]
rlabel metal2 19734 1622 19734 1622 0 wbs_sel_i[0]
rlabel metal2 21942 823 21942 823 0 wbs_sel_i[1]
rlabel metal2 24150 823 24150 823 0 wbs_sel_i[2]
rlabel metal2 26358 1044 26358 1044 0 wbs_sel_i[3]
rlabel metal2 16974 1588 16974 1588 0 wbs_stb_i
rlabel metal2 17526 1044 17526 1044 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 76000 87000
<< end >>
