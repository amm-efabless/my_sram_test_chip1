VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wishbone_sram
  CLASS BLOCK ;
  FOREIGN wishbone_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 380.000 BY 435.000 ;
  PIN sram_selected
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END sram_selected
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 9.180 5.200 10.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.180 5.200 60.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.180 5.200 110.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.180 5.200 160.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.180 5.200 210.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.180 5.200 260.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.180 5.200 310.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.180 5.200 360.940 430.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 9.560 375.140 11.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 59.560 375.140 61.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 109.560 375.140 111.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 159.560 375.140 161.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 209.560 375.140 211.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 259.560 375.140 261.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 309.560 375.140 311.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 359.560 375.140 361.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 409.560 375.140 411.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.510 0.000 11.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.510 0.000 41.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.510 0.000 71.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.510 0.000 101.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.510 0.000 131.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.510 0.000 161.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.510 0.000 191.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.510 0.000 221.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.510 0.000 251.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.510 0.000 281.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.510 0.000 311.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.510 0.000 341.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.510 0.000 371.610 435.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 20.940 5.200 22.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.940 5.200 72.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 120.940 5.200 122.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 170.940 5.200 172.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.940 5.200 222.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 270.940 5.200 272.700 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 320.940 5.200 322.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 370.940 5.200 372.700 430.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 21.320 375.140 23.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 71.320 375.140 73.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 121.320 375.140 123.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 171.320 375.140 173.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 221.320 375.140 223.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 271.320 375.140 273.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 321.320 375.140 323.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 371.320 375.140 373.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 421.320 375.140 423.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.510 0.000 26.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.510 0.000 56.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.510 0.000 86.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.510 0.000 116.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.510 0.000 146.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.510 0.000 176.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.510 0.000 206.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.510 0.000 236.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.510 0.000 266.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.510 0.000 296.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.510 0.000 326.610 435.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.510 0.000 356.610 435.000 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 374.900 429.845 ;
      LAYER met1 ;
        RECT 5.060 4.120 374.900 430.000 ;
      LAYER met2 ;
        RECT 10.100 30.140 358.900 427.870 ;
        RECT 10.100 30.000 20.660 30.140 ;
        RECT 11.220 4.920 20.660 30.000 ;
        RECT 22.980 4.920 58.900 30.140 ;
        RECT 61.220 4.920 70.660 30.140 ;
        RECT 72.980 4.920 108.900 30.140 ;
        RECT 111.220 4.920 120.660 30.140 ;
        RECT 122.980 4.920 158.900 30.140 ;
        RECT 161.220 4.920 170.660 30.140 ;
        RECT 172.980 4.920 208.900 30.140 ;
        RECT 211.220 4.920 220.660 30.140 ;
        RECT 222.980 4.920 258.900 30.140 ;
        RECT 261.220 30.000 308.900 30.140 ;
        RECT 261.220 4.920 270.660 30.000 ;
        RECT 272.980 4.920 308.900 30.000 ;
        RECT 311.220 4.920 320.660 30.140 ;
        RECT 322.980 4.920 358.900 30.140 ;
        RECT 361.220 4.920 366.520 427.870 ;
        RECT 10.100 4.280 366.520 4.920 ;
        RECT 10.100 3.670 15.450 4.280 ;
        RECT 16.290 3.670 73.410 4.280 ;
        RECT 74.250 3.670 76.170 4.280 ;
        RECT 77.010 3.670 78.930 4.280 ;
        RECT 79.770 3.670 81.690 4.280 ;
        RECT 82.530 3.670 84.450 4.280 ;
        RECT 85.290 3.670 87.210 4.280 ;
        RECT 88.050 3.670 89.970 4.280 ;
        RECT 90.810 3.670 92.730 4.280 ;
        RECT 93.570 3.670 95.490 4.280 ;
        RECT 96.330 3.670 98.250 4.280 ;
        RECT 99.090 3.670 101.010 4.280 ;
        RECT 101.850 3.670 103.770 4.280 ;
        RECT 104.610 3.670 106.530 4.280 ;
        RECT 107.370 3.670 109.290 4.280 ;
        RECT 110.130 3.670 112.050 4.280 ;
        RECT 112.890 3.670 114.810 4.280 ;
        RECT 115.650 3.670 117.570 4.280 ;
        RECT 118.410 3.670 120.330 4.280 ;
        RECT 121.170 3.670 123.090 4.280 ;
        RECT 123.930 3.670 125.850 4.280 ;
        RECT 126.690 3.670 128.610 4.280 ;
        RECT 129.450 3.670 131.370 4.280 ;
        RECT 132.210 3.670 134.130 4.280 ;
        RECT 134.970 3.670 136.890 4.280 ;
        RECT 137.730 3.670 139.650 4.280 ;
        RECT 140.490 3.670 142.410 4.280 ;
        RECT 143.250 3.670 145.170 4.280 ;
        RECT 146.010 3.670 147.930 4.280 ;
        RECT 148.770 3.670 150.690 4.280 ;
        RECT 151.530 3.670 153.450 4.280 ;
        RECT 154.290 3.670 156.210 4.280 ;
        RECT 157.050 3.670 158.970 4.280 ;
        RECT 159.810 3.670 161.730 4.280 ;
        RECT 162.570 3.670 164.490 4.280 ;
        RECT 165.330 3.670 167.250 4.280 ;
        RECT 168.090 3.670 170.010 4.280 ;
        RECT 170.850 3.670 172.770 4.280 ;
        RECT 173.610 3.670 175.530 4.280 ;
        RECT 176.370 3.670 178.290 4.280 ;
        RECT 179.130 3.670 181.050 4.280 ;
        RECT 181.890 3.670 183.810 4.280 ;
        RECT 184.650 3.670 186.570 4.280 ;
        RECT 187.410 3.670 189.330 4.280 ;
        RECT 190.170 3.670 192.090 4.280 ;
        RECT 192.930 3.670 194.850 4.280 ;
        RECT 195.690 3.670 197.610 4.280 ;
        RECT 198.450 3.670 200.370 4.280 ;
        RECT 201.210 3.670 203.130 4.280 ;
        RECT 203.970 3.670 205.890 4.280 ;
        RECT 206.730 3.670 208.650 4.280 ;
        RECT 209.490 3.670 211.410 4.280 ;
        RECT 212.250 3.670 214.170 4.280 ;
        RECT 215.010 3.670 216.930 4.280 ;
        RECT 217.770 3.670 219.690 4.280 ;
        RECT 220.530 3.670 222.450 4.280 ;
        RECT 223.290 3.670 225.210 4.280 ;
        RECT 226.050 3.670 227.970 4.280 ;
        RECT 228.810 3.670 230.730 4.280 ;
        RECT 231.570 3.670 233.490 4.280 ;
        RECT 234.330 3.670 236.250 4.280 ;
        RECT 237.090 3.670 239.010 4.280 ;
        RECT 239.850 3.670 241.770 4.280 ;
        RECT 242.610 3.670 244.530 4.280 ;
        RECT 245.370 3.670 247.290 4.280 ;
        RECT 248.130 3.670 250.050 4.280 ;
        RECT 250.890 3.670 252.810 4.280 ;
        RECT 253.650 3.670 255.570 4.280 ;
        RECT 256.410 3.670 258.330 4.280 ;
        RECT 259.170 3.670 261.090 4.280 ;
        RECT 261.930 3.670 263.850 4.280 ;
        RECT 264.690 3.670 266.610 4.280 ;
        RECT 267.450 3.670 269.370 4.280 ;
        RECT 270.210 3.670 272.130 4.280 ;
        RECT 272.970 3.670 274.890 4.280 ;
        RECT 275.730 3.670 277.650 4.280 ;
        RECT 278.490 3.670 280.410 4.280 ;
        RECT 281.250 3.670 283.170 4.280 ;
        RECT 284.010 3.670 285.930 4.280 ;
        RECT 286.770 3.670 288.690 4.280 ;
        RECT 289.530 3.670 291.450 4.280 ;
        RECT 292.290 3.670 294.210 4.280 ;
        RECT 295.050 3.670 296.970 4.280 ;
        RECT 297.810 3.670 299.730 4.280 ;
        RECT 300.570 3.670 302.490 4.280 ;
        RECT 303.330 3.670 305.250 4.280 ;
        RECT 306.090 3.670 308.010 4.280 ;
        RECT 308.850 3.670 310.770 4.280 ;
        RECT 311.610 3.670 313.530 4.280 ;
        RECT 314.370 3.670 316.290 4.280 ;
        RECT 317.130 3.670 319.050 4.280 ;
        RECT 319.890 3.670 321.810 4.280 ;
        RECT 322.650 3.670 324.570 4.280 ;
        RECT 325.410 3.670 327.330 4.280 ;
        RECT 328.170 3.670 330.090 4.280 ;
        RECT 330.930 3.670 332.850 4.280 ;
        RECT 333.690 3.670 335.610 4.280 ;
        RECT 336.450 3.670 338.370 4.280 ;
        RECT 339.210 3.670 341.130 4.280 ;
        RECT 341.970 3.670 343.890 4.280 ;
        RECT 344.730 3.670 346.650 4.280 ;
        RECT 347.490 3.670 349.410 4.280 ;
        RECT 350.250 3.670 352.170 4.280 ;
        RECT 353.010 3.670 354.930 4.280 ;
        RECT 355.770 3.670 357.690 4.280 ;
        RECT 358.530 3.670 360.450 4.280 ;
        RECT 361.290 3.670 363.210 4.280 ;
        RECT 364.050 3.670 366.520 4.280 ;
      LAYER met3 ;
        RECT 73.665 261.720 352.295 262.985 ;
        RECT 73.665 223.480 352.295 259.160 ;
        RECT 73.665 211.720 352.295 220.920 ;
        RECT 73.665 173.480 352.295 209.160 ;
        RECT 73.665 161.720 352.295 170.920 ;
        RECT 73.665 123.480 352.295 159.160 ;
        RECT 73.665 111.720 352.295 120.920 ;
        RECT 73.665 73.480 352.295 109.160 ;
        RECT 73.665 61.720 352.295 70.920 ;
        RECT 73.665 23.480 352.295 59.160 ;
        RECT 73.665 11.720 352.295 20.920 ;
        RECT 73.665 6.975 352.295 9.160 ;
      LAYER met4 ;
        RECT 199.935 16.495 203.110 262.985 ;
        RECT 207.010 16.495 218.110 262.985 ;
        RECT 222.010 16.495 233.110 262.985 ;
        RECT 237.010 16.495 248.110 262.985 ;
        RECT 252.010 16.495 263.110 262.985 ;
        RECT 267.010 16.495 278.110 262.985 ;
        RECT 282.010 16.495 293.110 262.985 ;
        RECT 297.010 16.495 308.110 262.985 ;
        RECT 312.010 16.495 323.110 262.985 ;
        RECT 327.010 16.495 338.110 262.985 ;
        RECT 342.010 16.495 342.865 262.985 ;
  END
END wishbone_sram
END LIBRARY

